magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1260 1520 1671
<< dnwell >>
rect 0 0 260 411
<< nwell >>
rect 0 0 260 411
<< nsubdiff >>
rect 0 368 260 375
rect 0 334 30 368
rect 64 334 113 368
rect 147 334 194 368
rect 228 334 260 368
rect 0 300 260 334
rect 0 266 30 300
rect 64 266 113 300
rect 147 266 194 300
rect 228 266 260 300
rect 0 232 260 266
rect 0 198 30 232
rect 64 198 113 232
rect 147 198 194 232
rect 228 198 260 232
rect 0 62 260 198
<< nsubdiffcont >>
rect 30 334 64 368
rect 113 334 147 368
rect 194 334 228 368
rect 30 266 64 300
rect 113 266 147 300
rect 194 266 228 300
rect 30 198 64 232
rect 113 198 147 232
rect 194 198 228 232
<< poly >>
rect 0 24 260 54
<< locali >>
rect 0 368 59 375
rect 93 368 260 375
rect 0 334 30 368
rect 93 341 113 368
rect 64 334 113 341
rect 147 334 194 368
rect 228 334 260 368
rect 0 303 260 334
rect 0 300 59 303
rect 93 300 260 303
rect 0 266 30 300
rect 93 269 113 300
rect 64 266 113 269
rect 147 266 194 300
rect 228 266 260 300
rect 0 232 260 266
rect 0 198 30 232
rect 64 198 113 232
rect 147 198 194 232
rect 228 198 260 232
rect 0 128 158 162
rect 192 128 260 162
rect 0 90 260 128
rect 0 56 158 90
rect 192 56 260 90
rect 0 55 260 56
rect 27 3 240 55
<< viali >>
rect 59 368 93 375
rect 59 341 64 368
rect 64 341 93 368
rect 59 300 93 303
rect 59 269 64 300
rect 64 269 93 300
rect 158 128 192 162
rect 158 56 192 90
<< metal1 >>
rect 0 219 18 411
rect 50 375 110 411
rect 50 341 59 375
rect 93 341 110 375
rect 50 303 110 341
rect 50 269 59 303
rect 93 269 110 303
rect 50 231 110 269
tri 50 220 61 231 ne
rect 61 220 110 231
tri 18 219 19 220 sw
tri 61 219 62 220 ne
rect 0 204 19 219
tri 19 204 34 219 sw
rect 0 146 34 204
rect 0 128 16 146
tri 16 128 34 146 nw
rect 0 0 14 128
tri 14 126 16 128 nw
tri 56 90 62 96 se
rect 62 90 110 220
tri 42 76 56 90 se
rect 56 76 110 90
rect 42 34 110 76
rect 42 0 76 34
tri 76 0 110 34 nw
rect 150 231 210 411
rect 150 221 200 231
tri 200 221 210 231 nw
rect 150 162 198 221
tri 198 219 200 221 nw
tri 240 219 242 221 se
rect 242 219 260 411
rect 150 128 158 162
rect 192 128 198 162
rect 150 90 198 128
tri 226 205 240 219 se
rect 240 205 260 219
rect 226 146 260 205
tri 226 126 246 146 ne
rect 150 56 158 90
rect 192 76 198 90
tri 198 76 218 96 sw
rect 192 56 218 76
rect 150 34 218 56
tri 150 0 184 34 ne
rect 184 0 218 34
rect 246 0 260 146
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_sp_colend_cent_ce.gds
string GDS_END 1954
string GDS_START 174
<< end >>
