# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_write_driver
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_write_driver ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.500000 BY  10.05500 ;
  PIN BL
    ANTENNADIFFAREA  0.270000 ;
    PORT
      LAYER met1 ;
        RECT 0.625000 9.505000 0.910000  9.795000 ;
        RECT 0.630000 9.795000 0.780000 10.055000 ;
    END
  END BL
  PIN BR
    ANTENNADIFFAREA  0.270000 ;
    PORT
      LAYER met1 ;
        RECT 1.510000 9.505000 1.795000  9.795000 ;
        RECT 1.640000 9.795000 1.790000 10.055000 ;
    END
  END BR
  PIN DIN
    ANTENNAGATEAREA  0.301500 ;
    PORT
      LAYER met1 ;
        RECT 1.275000 0.020000 1.575000 0.300000 ;
    END
  END DIN
  PIN E_N
    ANTENNAGATEAREA  0.330000 ;
    PORT
      LAYER met1 ;
        RECT 0.495000 0.470000 2.500000 0.640000 ;
        RECT 0.495000 0.640000 0.785000 0.780000 ;
    END
  END E_N
  PIN GND
    ANTENNADIFFAREA  0.177300 ;
    PORT
      LAYER met1 ;
        RECT 1.065000 7.775000 1.495000 7.805000 ;
        RECT 1.065000 7.805000 1.605000 7.975000 ;
        RECT 1.065000 7.975000 1.495000 8.005000 ;
      LAYER pwell ;
        RECT 1.145000 7.805000 1.605000 7.975000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.095000 2.920000 1.525000 3.150000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.670000 3.945000 2.100000 4.150000 ;
        RECT 1.735000 3.920000 2.100000 3.945000 ;
      LAYER pwell ;
        RECT 2.155000 3.640000 2.325000 4.100000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.386200 ;
    PORT
      LAYER met1 ;
        RECT 1.065000 5.590000 1.495000 5.820000 ;
      LAYER nwell ;
        RECT -0.760000 4.600000 3.280000 6.830000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.165000 0.840000 1.595000 1.070000 ;
      LAYER nwell ;
        RECT -0.760000 0.690000 3.280000 2.110000 ;
        RECT -0.760000 2.110000 3.270000 2.120000 ;
    END
  END VDD
  OBS
    LAYER li1 ;
      RECT 0.285000 5.570000 0.515000 5.900000 ;
      RECT 0.345000 0.870000 1.645000 1.040000 ;
      RECT 0.345000 1.040000 0.515000 1.880000 ;
      RECT 0.345000 2.050000 0.955000 2.220000 ;
      RECT 0.345000 2.220000 0.515000 5.570000 ;
      RECT 0.470000 0.500000 0.805000 0.670000 ;
      RECT 0.585000 7.900000 0.855000 8.235000 ;
      RECT 0.685000 3.650000 0.855000 4.420000 ;
      RECT 0.685000 4.420000 2.075000 4.590000 ;
      RECT 0.685000 4.590000 0.855000 5.350000 ;
      RECT 0.685000 6.080000 0.855000 7.900000 ;
      RECT 0.685000 8.545000 0.855000 9.735000 ;
      RECT 0.785000 1.290000 0.955000 2.050000 ;
      RECT 0.785000 2.440000 0.955000 3.030000 ;
      RECT 1.125000 4.760000 1.295000 5.620000 ;
      RECT 1.125000 5.620000 1.545000 5.790000 ;
      RECT 1.125000 5.790000 1.295000 6.665000 ;
      RECT 1.125000 7.165000 1.295000 7.805000 ;
      RECT 1.125000 7.805000 1.545000 7.975000 ;
      RECT 1.125000 7.975000 1.295000 9.635000 ;
      RECT 1.225000 0.840000 1.395000 0.870000 ;
      RECT 1.225000 1.040000 1.395000 1.880000 ;
      RECT 1.225000 2.440000 1.395000 3.120000 ;
      RECT 1.255000 0.100000 1.585000 0.270000 ;
      RECT 1.565000 3.660000 1.735000 3.950000 ;
      RECT 1.565000 3.950000 2.355000 4.120000 ;
      RECT 1.565000 4.120000 1.735000 4.250000 ;
      RECT 1.565000 4.590000 1.735000 5.350000 ;
      RECT 1.565000 6.080000 1.735000 6.825000 ;
      RECT 1.565000 6.825000 2.075000 6.995000 ;
      RECT 1.565000 6.995000 1.735000 7.565000 ;
      RECT 1.565000 8.545000 1.735000 9.735000 ;
      RECT 1.665000 1.290000 1.835000 1.950000 ;
      RECT 1.665000 1.950000 1.895000 2.120000 ;
      RECT 1.725000 2.120000 1.895000 2.890000 ;
      RECT 1.725000 2.890000 1.955000 2.990000 ;
      RECT 1.725000 2.990000 2.105000 3.110000 ;
      RECT 1.725000 3.110000 2.165000 3.160000 ;
      RECT 1.905000 4.590000 2.075000 5.570000 ;
      RECT 1.905000 5.570000 2.135000 5.900000 ;
      RECT 1.905000 6.995000 2.075000 9.615000 ;
      RECT 1.905000 9.615000 2.145000 9.945000 ;
      RECT 1.935000 3.160000 2.165000 3.490000 ;
      RECT 2.155000 3.700000 2.325000 3.950000 ;
    LAYER mcon ;
      RECT 0.555000 0.500000 0.725000 0.670000 ;
      RECT 0.685000 9.565000 0.855000 9.735000 ;
      RECT 1.225000 0.870000 1.395000 1.040000 ;
      RECT 1.225000 2.950000 1.395000 3.120000 ;
      RECT 1.335000 0.100000 1.505000 0.270000 ;
      RECT 1.565000 9.565000 1.735000 9.735000 ;
      RECT 1.800000 3.950000 1.970000 4.120000 ;
  END
END sky130_fd_bd_sram__openram_write_driver
END LIBRARY
