VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colend_cent_m2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colend_cent_m2 ;
  ORIGIN 0.055 -0.020 ;
  SIZE 1.410 BY 2.035 ;
  OBS
      LAYER met1 ;
        RECT 0.270 1.190 0.530 1.450 ;
        RECT -0.055 0.745 0.130 1.005 ;
        RECT 1.170 0.745 1.355 1.005 ;
        RECT 0.800 0.135 1.060 0.395 ;
      LAYER met2 ;
        RECT 0.000 1.600 1.300 2.055 ;
        RECT 0.000 1.180 1.300 1.460 ;
        RECT 0.000 1.005 1.300 1.030 ;
        RECT -0.055 0.745 1.355 1.005 ;
        RECT 0.000 0.580 1.300 0.745 ;
        RECT 0.000 0.020 1.300 0.405 ;
  END
END sky130_fd_bd_sram__sram_sp_colend_cent_m2
END LIBRARY

