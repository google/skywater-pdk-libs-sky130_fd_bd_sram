magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1246 -1260 1500 1279
<< locali >>
rect 14 0 240 19
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_colend_half_limcon_opta.gds
string GDS_END 258
string GDS_START 190
<< end >>
