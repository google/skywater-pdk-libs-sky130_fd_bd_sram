# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_nand2_dec
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_nand2_dec ;
  ORIGIN -0.290000 -0.265000 ;
  SIZE  4.285000 BY  1.715000 ;
  PIN GND
    ANTENNADIFFAREA  0.297600 ;
    PORT
      LAYER met1 ;
        RECT 0.380000 0.440000 0.620000 0.500000 ;
        RECT 0.380000 0.500000 1.470000 0.680000 ;
        RECT 0.380000 0.680000 0.620000 0.740000 ;
        RECT 1.230000 0.145000 1.470000 0.500000 ;
        RECT 1.230000 0.680000 1.470000 2.010000 ;
      LAYER pwell ;
        RECT 0.290000 0.500000 0.710000 0.680000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.415800 ;
    PORT
      LAYER met1 ;
        RECT 3.350000 0.150000 3.600000 0.680000 ;
        RECT 3.350000 0.680000 4.560000 0.850000 ;
        RECT 3.350000 0.850000 3.600000 2.010000 ;
        RECT 4.225000 0.850000 4.560000 0.890000 ;
        RECT 4.245000 0.640000 4.560000 0.680000 ;
      LAYER nwell ;
        RECT 2.060000 -0.300000 4.880000 2.390000 ;
    END
  END VDD
  OBS
    LAYER li1 ;
      RECT 0.330000 0.500000 0.710000 0.680000 ;
      RECT 0.350000 0.870000 0.680000 1.040000 ;
      RECT 0.350000 1.410000 0.680000 1.580000 ;
      RECT 1.040000 0.710000 1.700000 0.880000 ;
      RECT 1.050000 1.570000 4.440000 1.740000 ;
      RECT 2.545000 0.670000 2.860000 0.675000 ;
      RECT 2.545000 0.675000 3.425000 0.680000 ;
      RECT 2.545000 0.680000 3.640000 0.845000 ;
      RECT 2.545000 0.845000 2.990000 0.850000 ;
      RECT 2.545000 0.850000 2.715000 1.570000 ;
      RECT 3.300000 0.845000 3.640000 0.850000 ;
      RECT 3.300000 1.130000 3.635000 1.300000 ;
      RECT 4.225000 0.680000 4.575000 0.860000 ;
    LAYER mcon ;
      RECT 0.415000 0.505000 0.585000 0.675000 ;
      RECT 1.270000 0.710000 1.440000 0.880000 ;
      RECT 3.385000 1.130000 3.555000 1.300000 ;
      RECT 4.315000 0.685000 4.485000 0.855000 ;
  END
END sky130_fd_bd_sram__openram_nand2_dec
END LIBRARY
