# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_cell_1rw_1r_cap_row
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_cell_1rw_1r_cap_row ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.120000 BY  1.975000 ;
  OBS
    LAYER met2 ;
      RECT -0.210000 -0.275000 3.120000 0.275000 ;
      RECT -0.210000  0.515000 3.120000 0.755000 ;
      RECT -0.210000  0.995000 2.020000 1.065000 ;
      RECT -0.210000  1.065000 3.120000 1.305000 ;
      RECT -0.210000  1.305000 2.020000 1.375000 ;
      RECT -0.210000  1.615000 3.120000 1.855000 ;
      RECT  2.190000  0.755000 2.600000 0.825000 ;
      RECT  2.190000  1.545000 2.600000 1.615000 ;
      RECT  2.770000  0.995000 3.120000 1.065000 ;
      RECT  2.770000  1.305000 3.120000 1.375000 ;
  END
END sky130_fd_bd_sram__openram_cell_1rw_1r_cap_row
END LIBRARY
