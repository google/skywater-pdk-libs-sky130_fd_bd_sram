magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1295 -1260 1338 1576
<< metal1 >>
rect 0 180 78 316
rect -35 128 78 180
rect 42 0 78 128
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_swldrv_strap1.gds
string GDS_END 270
string GDS_START 170
<< end >>
