* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_metopt1.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_metopt1
.ends
