# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_met23_1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_met23_1 ;
  ORIGIN  3.110000  0.055000 ;
  SIZE  3.165000 BY  1.690000 ;
  OBS
    LAYER met1 ;
      RECT -3.110000  1.450000 -2.925000 1.635000 ;
      RECT -0.130000 -0.055000  0.055000 0.130000 ;
      RECT -0.130000  1.450000  0.055000 1.635000 ;
    LAYER met2 ;
      RECT -3.110000  1.450000 -2.815000 1.580000 ;
      RECT -3.110000  1.580000 -2.915000 1.620000 ;
      RECT -3.110000  1.620000 -2.925000 1.635000 ;
      RECT -3.095000  1.440000 -2.815000 1.450000 ;
      RECT -3.055000  0.675000 -0.975000 1.100000 ;
      RECT -3.055000  1.340000 -2.815000 1.440000 ;
      RECT -2.840000  0.000000 -2.360000 0.240000 ;
      RECT -2.740000 -0.040000 -2.460000 0.000000 ;
      RECT -1.455000  0.000000  0.055000 0.130000 ;
      RECT -1.455000  0.130000  0.000000 0.185000 ;
      RECT -1.455000  0.185000 -0.975000 0.675000 ;
      RECT -1.455000  1.100000 -0.975000 1.395000 ;
      RECT -1.455000  1.395000  0.000000 1.450000 ;
      RECT -1.455000  1.450000  0.055000 1.580000 ;
      RECT -0.130000 -0.055000  0.055000 0.000000 ;
      RECT -0.130000  1.580000  0.055000 1.635000 ;
    LAYER met3 ;
      RECT -3.095000  1.440000  0.000000 1.580000 ;
      RECT -3.095000  1.580000 -2.915000 1.620000 ;
      RECT -3.055000  0.000000  0.000000 0.205000 ;
      RECT -3.055000  0.505000  0.000000 1.075000 ;
      RECT -3.055000  1.375000  0.000000 1.440000 ;
      RECT -2.740000 -0.040000 -2.460000 0.000000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_met23_1
END LIBRARY
