* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_ce.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_ce
X0 a_174_0# a_0_24# a_174_0# w_96_0# sky130_fd_pr__nfet_01v8 ad=1.68e+10p pd=520000u as=0p ps=0u w=70000u l=210000u
.ends
