magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1201 1500 1517
<< metal2 >>
rect 0 213 240 257
rect 191 205 240 213
rect 0 171 58 179
rect 0 127 240 171
rect 0 59 240 93
<< properties >>
string GDS_FILE sky130_fd_bd_sram__openram_sp_cell_met2.gds
string GDS_END 398
string GDS_START 170
<< end >>
