VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell_p1_serif
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell_p1_serif ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END sky130_fd_bd_sram__sram_sp_cell_p1_serif
END LIBRARY

