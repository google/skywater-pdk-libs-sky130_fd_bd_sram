# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_tap
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_tap ;
  ORIGIN  0.000000  0.310000 ;
  SIZE  2.595000 BY  0.545000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.310000 0.165000 -0.150000 ;
      RECT 0.000000 -0.150000 1.180000  0.150000 ;
      RECT 0.000000  0.150000 1.310000  0.235000 ;
    LAYER pwell ;
      RECT 0.000000 -0.140000 1.510000 0.075000 ;
      RECT 0.000000  0.075000 1.575000 0.235000 ;
      RECT 2.095000  0.035000 2.595000 0.235000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_tap
END LIBRARY
