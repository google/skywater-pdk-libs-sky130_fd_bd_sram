magic
tech sky130A
magscale 1 2
timestamp 1621288227
<< dnwell >>
rect 0 0 260 411
<< nwell >>
rect 0 0 260 411
<< nsubdiff >>
rect 0 368 260 375
rect 0 334 30 368
rect 64 334 113 368
rect 147 334 194 368
rect 228 334 260 368
rect 0 300 260 334
rect 0 266 30 300
rect 64 266 113 300
rect 147 266 194 300
rect 228 266 260 300
rect 0 232 260 266
rect 0 198 30 232
rect 64 198 113 232
rect 147 198 194 232
rect 228 198 260 232
rect 0 62 260 198
<< nsubdiffcont >>
rect 30 334 64 368
rect 113 334 147 368
rect 194 334 228 368
rect 30 266 64 300
rect 113 266 147 300
rect 194 266 228 300
rect 30 198 64 232
rect 113 198 147 232
rect 194 198 228 232
<< poly >>
rect 0 24 260 54
<< locali >>
rect 0 368 59 375
rect 93 368 260 375
rect 0 334 30 368
rect 93 341 113 368
rect 64 334 113 341
rect 147 334 194 368
rect 228 334 260 368
rect 0 303 260 334
rect 0 300 59 303
rect 93 300 260 303
rect 0 266 30 300
rect 93 269 113 300
rect 64 266 113 269
rect 147 266 194 300
rect 228 266 260 300
rect 0 232 260 266
rect 0 198 30 232
rect 64 198 113 232
rect 147 198 194 232
rect 228 198 260 232
rect 0 128 158 162
rect 192 128 260 162
rect 0 90 260 128
rect 0 56 158 90
rect 192 56 260 90
rect 0 55 260 56
rect 27 3 240 55
<< viali >>
rect 59 368 93 375
rect 59 341 64 368
rect 64 341 93 368
rect 59 300 93 303
rect 59 269 64 300
rect 64 269 93 300
rect 158 128 192 162
rect 158 56 192 90
<< metal1 >>
rect 0 204 18 411
rect 50 375 110 411
rect 50 341 59 375
rect 93 341 110 375
rect 50 303 110 341
rect 50 289 59 303
rect 93 289 110 303
rect 50 239 55 289
rect 105 239 110 289
rect 50 231 110 239
tri 18 204 34 220 sw
tri 50 219 62 231 ne
rect 0 200 34 204
rect 25 150 34 200
rect 0 146 34 150
rect 0 0 14 146
tri 14 126 34 146 nw
tri 42 76 62 96 se
rect 62 76 110 231
rect 42 34 110 76
rect 42 0 76 34
tri 76 0 110 34 nw
rect 150 231 210 411
rect 150 162 198 231
tri 198 219 210 231 nw
rect 150 128 158 162
rect 192 128 198 162
rect 150 90 198 128
tri 226 205 242 221 se
rect 242 205 260 411
rect 226 200 260 205
rect 226 150 235 200
rect 226 146 260 150
tri 226 126 246 146 ne
rect 150 56 158 90
rect 192 78 198 90
tri 198 78 216 96 sw
rect 211 76 216 78
tri 216 76 218 78 sw
rect 150 34 161 56
tri 150 28 156 34 ne
rect 156 28 161 34
rect 211 28 218 76
tri 156 0 184 28 ne
rect 184 0 218 28
rect 246 0 260 146
<< via1 >>
rect 55 269 59 289
rect 59 269 93 289
rect 93 269 105 289
rect 55 239 105 269
rect -10 150 25 200
rect 235 150 270 200
rect 161 56 192 78
rect 192 56 211 78
rect 161 28 211 56
<< metal2 >>
rect 0 320 260 411
rect 0 289 260 292
rect 0 239 55 289
rect 105 239 260 289
rect 0 236 260 239
rect 0 200 260 206
rect 25 150 235 200
rect 0 116 260 150
rect 0 78 260 81
rect 0 28 161 78
rect 211 28 260 78
rect 0 4 260 28
<< labels >>
rlabel metal1 s 246 0 260 19 4 VPWR
rlabel metal1 s 154 162 198 198 4 VNB
rlabel metal1 s 62 162 106 198 4 VPB
rlabel metal1 s 0 0 14 19 4 VPWR
<< end >>
