# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_cell_6t
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_cell_6t ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.500000 BY  1.580000 ;
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.660000 0.170000 0.710000 0.230000 ;
    END
  END VNB
  PIN VPB
    ANTENNADIFFAREA  0.442800 ;
    PORT
      LAYER met2 ;
        RECT -0.650000 1.065000 3.150000 1.285000 ;
        RECT  1.605000 1.025000 3.150000 1.065000 ;
      LAYER nwell ;
        RECT 1.340000 0.065000 3.150000 1.515000 ;
        RECT 1.370000 0.000000 3.150000 0.065000 ;
        RECT 1.370000 1.515000 3.150000 1.580000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      POLYGON  0.955000  1.150000  1.005000 1.150000 0.955000 1.100000 ;
      POLYGON  1.580000  0.475000  1.580000 0.415000 1.520000 0.415000 ;
      RECT -0.370000  0.200000 -0.200000 0.370000 ;
      RECT -0.085000  0.160000  0.085000 0.330000 ;
      RECT -0.085000  0.715000  0.085000 0.885000 ;
      RECT -0.085000  1.055000  0.085000 1.225000 ;
      RECT  0.175000  0.605000  0.345000 0.775000 ;
      RECT  0.175000  0.965000  0.345000 1.135000 ;
      RECT  0.200000  0.200000  0.370000 0.370000 ;
      RECT  0.565000  0.705000  0.735000 0.875000 ;
      RECT  0.840000 -0.075000  0.980000 0.075000 ;
      RECT  0.840000  0.310000  0.980000 0.395000 ;
      RECT  0.840000  0.395000  1.000000 0.480000 ;
      RECT  0.840000  1.100000  0.955000 1.150000 ;
      RECT  0.840000  1.150000  1.005000 1.185000 ;
      RECT  0.840000  1.185000  0.980000 1.270000 ;
      RECT  0.840000  1.505000  0.980000 1.655000 ;
      RECT  0.985000  1.495000  1.155000 1.665000 ;
      RECT  1.185000  0.520000  1.355000 0.670000 ;
      RECT  1.185000  0.910000  1.355000 1.060000 ;
      RECT  1.345000 -0.085000  1.515000 0.085000 ;
      RECT  1.520000  0.305000  1.660000 0.415000 ;
      RECT  1.520000  1.105000  1.660000 1.275000 ;
      RECT  1.580000  0.415000  1.660000 0.475000 ;
      RECT  1.765000  0.705000  1.935000 0.875000 ;
      RECT  2.155000  0.605000  2.325000 0.775000 ;
      RECT  2.155000  0.965000  2.325000 1.135000 ;
      RECT  2.245000  0.200000  2.755000 0.370000 ;
      RECT  2.415000  0.620000  2.585000 0.790000 ;
      RECT  2.415000  0.960000  2.585000 1.130000 ;
    LAYER mcon ;
      RECT 2.415000 0.200000 2.585000 0.370000 ;
    LAYER met1 ;
      POLYGON -0.130000  0.105000 -0.095000 0.105000 -0.095000 0.070000 ;
      POLYGON -0.095000  0.410000 -0.095000 0.375000 -0.130000 0.375000 ;
      POLYGON  0.095000  0.105000  0.130000 0.105000  0.095000 0.070000 ;
      POLYGON  0.095000  0.410000  0.130000 0.375000  0.095000 0.375000 ;
      POLYGON  0.140000  0.580000  0.270000 0.580000  0.270000 0.450000 ;
      POLYGON  0.380000  0.570000  0.440000 0.510000  0.380000 0.510000 ;
      POLYGON  0.520000  0.630000  0.545000 0.630000  0.545000 0.605000 ;
      POLYGON  1.735000  0.645000  1.745000 0.645000  1.745000 0.635000 ;
      POLYGON  1.955000  0.645000  1.965000 0.645000  1.955000 0.635000 ;
      POLYGON  2.120000  0.600000  2.120000 0.540000  2.060000 0.540000 ;
      POLYGON  2.230000  0.600000  2.350000 0.600000  2.230000 0.480000 ;
      POLYGON  2.350000  0.610000  2.360000 0.610000  2.350000 0.600000 ;
      POLYGON  2.370000  0.100000  2.400000 0.100000  2.400000 0.070000 ;
      POLYGON  2.390000  0.440000  2.390000 0.420000  2.370000 0.420000 ;
      POLYGON  2.600000  0.100000  2.630000 0.100000  2.600000 0.070000 ;
      POLYGON  2.610000  0.440000  2.630000 0.420000  2.610000 0.420000 ;
      RECT -0.130000  0.105000  0.130000 0.375000 ;
      RECT -0.095000  0.070000  0.095000 0.105000 ;
      RECT -0.095000  0.375000  0.095000 0.410000 ;
      RECT  0.000000  0.795000  0.780000 0.925000 ;
      RECT  0.000000  0.925000  0.720000 1.035000 ;
      RECT  0.140000  0.580000  0.380000 0.795000 ;
      RECT  0.140000  1.035000  0.380000 1.580000 ;
      RECT  0.270000  0.000000  0.440000 0.510000 ;
      RECT  0.270000  0.510000  0.380000 0.580000 ;
      RECT  0.520000  0.630000  0.780000 0.795000 ;
      RECT  0.520000  1.035000  0.720000 1.315000 ;
      RECT  0.545000  0.605000  0.780000 0.630000 ;
      RECT  0.580000 -0.075000  0.720000 0.605000 ;
      RECT  0.580000  1.315000  0.720000 1.580000 ;
      RECT  0.950000  1.435000  1.190000 1.725000 ;
      RECT  1.000000  0.000000  1.140000 1.435000 ;
      RECT  1.310000 -0.145000  1.550000 0.145000 ;
      RECT  1.360000  0.145000  1.500000 1.580000 ;
      RECT  1.720000  0.990000  2.500000 1.035000 ;
      RECT  1.720000  1.035000  1.980000 1.315000 ;
      RECT  1.735000  0.645000  1.965000 0.795000 ;
      RECT  1.735000  0.795000  2.500000 0.990000 ;
      RECT  1.745000  0.635000  1.955000 0.645000 ;
      RECT  1.780000 -0.075000  1.920000 0.635000 ;
      RECT  1.780000  1.315000  1.920000 1.580000 ;
      RECT  2.060000  0.000000  2.230000 0.540000 ;
      RECT  2.120000  0.540000  2.230000 0.600000 ;
      RECT  2.120000  0.600000  2.350000 0.610000 ;
      RECT  2.120000  0.610000  2.360000 0.795000 ;
      RECT  2.120000  1.035000  2.360000 1.580000 ;
      RECT  2.370000  0.100000  2.630000 0.420000 ;
      RECT  2.390000  0.420000  2.610000 0.440000 ;
      RECT  2.400000  0.070000  2.600000 0.100000 ;
    LAYER met2 ;
      RECT -0.650000 0.295000 3.150000 0.465000 ;
      RECT -0.650000 0.635000 3.150000 0.855000 ;
      RECT -0.650000 0.855000 0.940000 0.895000 ;
      RECT -0.160000 0.120000 0.160000 0.295000 ;
      RECT -0.130000 0.115000 0.130000 0.120000 ;
      RECT  2.370000 0.120000 2.630000 0.295000 ;
    LAYER pwell ;
      RECT -0.235000 0.610000 0.235000 1.260000 ;
    LAYER via ;
      RECT -0.130000 0.115000 0.130000 0.375000 ;
      RECT  0.520000 0.635000 0.780000 0.895000 ;
      RECT  1.720000 1.025000 1.980000 1.285000 ;
      RECT  2.370000 0.150000 2.630000 0.410000 ;
  END
END sky130_fd_bd_sram__openram_cell_6t
END LIBRARY
