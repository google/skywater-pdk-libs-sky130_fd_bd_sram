* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda_p1m_siz.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda_p1m_siz
.ends
