# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_horstrap_half
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_horstrap_half ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.200000 BY  0.790000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.305000 1.200000 0.485000 ;
    LAYER mcon ;
      RECT 0.000000 0.310000 0.085000 0.480000 ;
    LAYER met1 ;
      RECT 0.000000 0.205000 0.210000 0.585000 ;
      RECT 0.390000 0.000000 0.570000 0.790000 ;
      RECT 0.750000 0.000000 0.930000 0.790000 ;
      RECT 1.110000 0.000000 1.200000 0.790000 ;
    LAYER met2 ;
      RECT 0.000000 0.120000 1.200000 0.670000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 1.200000 0.205000 ;
      RECT 0.000000 0.585000 1.200000 0.790000 ;
    LAYER nwell ;
      RECT 0.720000 0.000000 1.200000 0.790000 ;
    LAYER pwell ;
      RECT 0.190000 0.200000 0.400000 0.590000 ;
  END
END sky130_fd_bd_sram__sram_dp_horstrap_half
END LIBRARY
