magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1271 1882 1429
<< via1 >>
rect -11 132 26 169
rect 585 132 622 169
rect -11 -11 26 26
rect 585 -11 622 26
<< metal2 >>
rect 28 130 48 158
rect 0 28 48 130
rect 28 0 48 28
rect 320 132 585 158
rect 320 26 611 132
rect 320 0 585 26
<< via2 >>
rect -8 132 26 166
rect 26 132 28 166
rect -8 130 28 132
rect -8 26 28 28
rect -8 -8 26 26
rect 26 -8 28 26
<< metal3 >>
rect 28 130 611 158
rect 0 117 611 130
rect 0 41 41 117
rect 0 28 611 41
rect 28 0 611 28
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_blkinv_met23.gds
string GDS_END 878
string GDS_START 170
<< end >>
