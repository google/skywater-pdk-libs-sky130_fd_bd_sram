* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__sram_dp_swldrv_base a_n70_24# m1_n403_0# m1_n223_0# SUBS
+ a_n287_182# w_n611_0# a_n517_117# w_n192_0# a_n517_27#
X0 a_n517_117# a_n611_0# a_n517_27# w_n611_0# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 SUBS a_n287_182# a_n517_117# SUBS sky130_fd_pr__nfet_01v8 w=500000u l=150000u
X2 a_n517_117# a_n611_0# SUBS SUBS sky130_fd_pr__nfet_01v8 w=500000u l=150000u
.ends
* Top level circuit sky130_fd_bd_sram__sram_dp_swldrv_opt1a
Xsky130_fd_bd_sram__sram_dp_swldrv_base_0 a_567_24# sky130_fd_bd_sram__sram_dp_swldrv_mcon_0/li_0_14#
+ sky130_fd_bd_sram__sram_dp_swldrv_base_0/m1_n223_0# SUBS sky130_fd_bd_sram__sram_dp_swldrv_base_0/m1_n223_0#
+ sky130_fd_bd_sram__sram_dp_swldrv_tap_0/a_0_n28# a_567_24# SUBS sky130_fd_bd_sram__sram_dp_swldrv_mcon_0/li_0_14#
+ sky130_fd_bd_sram__sram_dp_swldrv_base
.end
