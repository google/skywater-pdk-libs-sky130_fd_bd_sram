magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1263 1872 1454
<< nwell >>
rect 64 158 322 194
rect 0 0 351 158
<< nmos >>
rect 419 116 481 146
rect 419 12 481 42
<< pmos >>
rect 100 128 286 158
rect 100 42 286 72
<< ndiff >>
rect 419 146 481 158
rect 419 96 481 116
rect 419 62 431 96
rect 465 62 481 96
rect 419 42 481 62
rect 419 0 481 12
<< pdiff >>
rect 100 158 286 159
rect 100 117 286 128
rect 100 83 172 117
rect 206 83 240 117
rect 274 83 286 117
rect 100 72 286 83
rect 100 31 286 42
rect 100 0 118 31
rect 152 0 210 31
rect 244 0 286 31
<< ndiffc >>
rect 431 62 465 96
<< pdiffc >>
rect 172 83 206 117
rect 240 83 274 117
rect 118 0 152 31
rect 210 0 244 31
<< poly >>
rect 48 128 100 158
rect 286 128 312 158
rect 48 72 78 128
rect 365 116 419 146
rect 481 116 509 146
rect 365 72 395 116
rect 48 42 100 72
rect 286 42 395 72
rect 559 104 611 134
rect 559 96 609 104
rect 559 62 567 96
rect 601 62 609 96
rect 559 54 609 62
rect 365 12 419 42
rect 481 12 509 42
rect 559 24 611 54
<< polycont >>
rect 567 62 601 96
<< locali >>
rect 102 31 136 158
rect 459 141 493 158
rect 527 141 576 148
rect 172 117 222 133
rect 459 124 576 141
rect 499 120 576 124
rect 206 83 240 117
rect 274 106 330 117
rect 274 83 431 106
rect 517 105 576 120
rect 517 96 611 105
rect 172 67 431 83
rect 296 52 431 67
rect 465 62 481 96
rect 517 62 567 96
rect 517 53 611 62
rect 517 38 576 53
rect 499 34 576 38
rect 102 0 118 31
rect 152 0 210 31
rect 244 0 260 31
rect 459 17 576 34
rect 459 0 493 17
rect 527 10 576 17
rect 102 -3 260 0
<< viali >>
rect 493 141 527 158
rect 594 62 601 96
rect 601 62 611 96
rect 493 0 527 17
<< metal1 >>
rect 0 0 78 158
rect 118 0 168 158
rect 208 0 258 158
rect 298 0 348 158
rect 388 0 438 158
rect 487 141 493 158
rect 527 141 611 158
rect 487 96 611 141
rect 487 62 594 96
rect 487 17 611 62
rect 487 0 493 17
rect 527 0 611 17
use sky130_fd_bd_sram__sram_dp_blkinv_p1m_siz  sky130_fd_bd_sram__sram_dp_blkinv_p1m_siz_0
timestamp 0
transform 1 0 90 0 1 18
box 469 6 470 117
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_0
timestamp 0
transform 1 0 257 0 1 100
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_1
timestamp 0
transform 1 0 189 0 1 100
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_2
timestamp 0
transform 1 0 135 0 1 14
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_3
timestamp 0
transform 1 0 227 0 1 14
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_4
timestamp 0
transform 1 0 448 0 1 79
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_licon_1  sky130_fd_bd_sram__sram_dp_licon_1_5
timestamp 0
transform 1 0 584 0 1 79
box 0 -1 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_li_drop  sky130_fd_bd_sram__sram_dp_swldrv_li_drop_0
timestamp 0
transform 1 0 611 0 1 0
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_li_drop  sky130_fd_bd_sram__sram_dp_swldrv_li_drop_1
timestamp 0
transform 1 0 611 0 -1 158
box 0 0 1 1
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_blkinv_base.gds
string GDS_END 4066
string GDS_START 1558
<< end >>
