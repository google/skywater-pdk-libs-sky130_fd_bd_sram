# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_mcon
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_mcon ;
  ORIGIN  0.045000  0.020000 ;
  SIZE  1.160000 BY  1.360000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.070000 0.170000 0.240000 ;
      RECT 0.900000 1.080000 1.070000 1.250000 ;
    LAYER met1 ;
      RECT -0.045000 -0.020000 0.215000 0.330000 ;
      RECT  0.855000  0.990000 1.115000 1.340000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_mcon
END LIBRARY
