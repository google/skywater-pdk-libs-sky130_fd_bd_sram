VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colend_p_cent_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colend_p_cent_ce ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.300 BY 2.055 ;
  OBS
      LAYER pwell ;
        RECT 0.000 0.530 1.300 1.680 ;
      LAYER li1 ;
        RECT 0.000 1.175 1.300 1.875 ;
        RECT 0.000 0.275 1.300 1.005 ;
        RECT 0.135 0.015 1.200 0.275 ;
      LAYER mcon ;
        RECT 0.350 1.705 0.520 1.875 ;
        RECT 0.350 1.345 0.520 1.515 ;
        RECT 0.790 0.640 0.960 0.810 ;
        RECT 0.790 0.280 0.960 0.450 ;
      LAYER met1 ;
        RECT 0.000 1.685 0.150 2.055 ;
        RECT 0.000 1.020 0.090 1.685 ;
        POLYGON 0.090 1.685 0.150 1.685 0.090 1.625 ;
        POLYGON 0.310 1.615 0.310 1.555 0.250 1.555 ;
        RECT 0.310 1.555 0.550 2.055 ;
        RECT 0.250 1.155 0.550 1.555 ;
        POLYGON 0.250 1.155 0.305 1.155 0.305 1.100 ;
        RECT 0.305 1.100 0.550 1.155 ;
        POLYGON 0.090 1.100 0.170 1.020 0.090 1.020 ;
        POLYGON 0.305 1.100 0.310 1.100 0.310 1.095 ;
        RECT 0.000 0.730 0.170 1.020 ;
        RECT 0.000 0.000 0.070 0.730 ;
        POLYGON 0.070 0.730 0.170 0.730 0.070 0.630 ;
        POLYGON 0.310 0.480 0.310 0.380 0.210 0.380 ;
        RECT 0.310 0.380 0.550 1.100 ;
        RECT 0.210 0.170 0.550 0.380 ;
        RECT 0.210 0.000 0.380 0.170 ;
        POLYGON 0.380 0.170 0.550 0.170 0.380 0.000 ;
        RECT 0.750 1.555 0.990 2.055 ;
        RECT 1.150 1.685 1.300 2.055 ;
        POLYGON 1.150 1.685 1.210 1.685 1.210 1.625 ;
        POLYGON 0.990 1.615 1.050 1.555 0.990 1.555 ;
        RECT 0.750 1.155 1.050 1.555 ;
        RECT 0.750 0.380 0.990 1.155 ;
        POLYGON 0.990 1.155 1.050 1.155 0.990 1.095 ;
        POLYGON 1.210 1.105 1.210 1.095 1.200 1.095 ;
        RECT 1.210 1.095 1.300 1.685 ;
        POLYGON 1.200 1.095 1.200 1.025 1.130 1.025 ;
        RECT 1.200 1.025 1.300 1.095 ;
        RECT 1.130 0.730 1.300 1.025 ;
        POLYGON 1.130 0.730 1.230 0.730 1.230 0.630 ;
        POLYGON 0.990 0.480 1.090 0.380 0.990 0.380 ;
        RECT 0.750 0.170 1.090 0.380 ;
        POLYGON 0.750 0.170 0.920 0.170 0.920 0.000 ;
        RECT 0.920 0.000 1.090 0.170 ;
        RECT 1.230 0.000 1.300 0.730 ;
  END
END sky130_fd_bd_sram__sram_sp_colend_p_cent_ce
END LIBRARY

