# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_strap2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_strap2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.370000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT 0.050000 0.155000 0.220000 0.325000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 0.370000 0.440000 ;
      RECT 0.000000 0.900000 0.185000 1.580000 ;
    LAYER met2 ;
      RECT 0.025000 0.000000 0.345000 0.435000 ;
    LAYER via ;
      RECT 0.055000 0.100000 0.315000 0.360000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_strap2
END LIBRARY
