
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.SUBCKT sky130_fd_bd_sram__openram_cell_6t bl br wl vdd gnd
* Inverter 1
Mnpd_bar Qbar Q gnd gnd npd W=0.210 L=0.150 m=1 mult=1
Mppu_bar Qbar Q vdd vdd pp W=0.140 L=0.150 m=1 mult=1

* Inverer 2
Mnpd_tr Q Qbar gnd gnd npd W=0.210 L=0.150 m=1 mult=1
Mppu_tr Q Qbar vdd vdd pp W=0.140 L=0.150 m=1 mult=1

* Access transistors
Mspecial_nfet_pass_tr bl wl Q gnd special_nfet_pass W=0.140 L=0.150 m=1 mult=1
Mspecial_nfet_pass_bar br wl Qbar gnd special_nfet_pass W=0.140 L=0.150 m=1 mult=1

* Parasitic transistors
Mpdo_tr Q wl Q vdd pp W=0.140 L=0.25 m=1 mult=1
Mpdo_bar Qbar wl Qbar vdd pp W=0.140 L=0.25 m=1 mult=1

.ENDS sky130_fd_bd_sram__openram_cell_6t
