magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1390 -1289 1890 1605
<< dnwell >>
rect -130 0 630 316
<< nwell >>
rect 274 303 630 316
rect 268 13 630 303
rect 274 0 630 13
<< pwell >>
rect -47 122 47 252
rect 132 34 142 46
<< npd >>
rect 168 262 196 292
rect 168 182 210 212
rect 168 104 210 134
rect 168 24 196 54
<< pmoshvt >>
rect 304 262 332 267
rect 304 182 332 212
rect 304 104 332 134
rect 304 49 332 54
<< ndiff >>
rect 168 292 196 301
rect 168 254 196 262
tri 191 220 201 230 se
rect 201 220 210 237
rect 168 212 210 220
rect 168 174 210 182
rect 103 142 116 174
rect 144 142 210 174
rect 168 134 210 142
rect 168 96 210 104
rect 200 79 210 96
rect 168 54 196 62
rect 168 15 196 24
<< pdiff >>
rect 304 255 332 262
rect 304 212 332 221
rect 304 174 332 182
rect 304 142 356 174
rect 384 142 397 174
rect 304 134 332 142
rect 304 95 332 104
tri 304 83 316 95 nw
rect 304 54 332 61
<< ndiffc >>
rect 168 301 196 331
rect 168 237 196 254
rect 168 230 201 237
rect 168 220 191 230
tri 191 220 201 230 nw
rect 116 142 144 174
rect 168 79 200 96
rect 168 62 196 79
rect 168 -15 196 15
<< pdiffc >>
rect 304 221 332 255
rect 356 142 384 174
tri 304 83 316 95 se
rect 316 83 332 95
rect 304 61 332 83
<< psubdiff >>
rect -47 245 47 252
rect -47 211 -17 245
rect 17 211 47 245
rect -47 177 47 211
rect -47 143 -17 177
rect 17 143 47 177
rect -47 122 47 143
<< nsubdiff >>
rect 453 226 547 252
rect 453 192 483 226
rect 517 192 547 226
rect 453 158 547 192
rect 453 124 483 158
rect 517 124 547 158
rect 453 100 547 124
<< psubdiffcont >>
rect -17 211 17 245
rect -17 143 17 177
<< nsubdiffcont >>
rect 483 192 517 226
rect 483 124 517 158
<< poly >>
rect -130 262 168 292
rect 196 267 630 292
rect 196 262 304 267
rect 332 262 630 267
rect -90 90 -57 262
rect 57 90 90 262
rect 146 182 168 212
rect 210 182 237 212
rect 271 182 304 212
rect 332 182 354 212
rect 146 104 168 134
rect 210 104 237 134
rect 271 104 304 134
rect 332 104 354 134
rect -90 74 90 90
rect -90 54 -74 74
rect -130 40 -74 54
rect -40 40 40 74
rect 74 54 90 74
rect 410 90 443 262
rect 557 90 590 262
rect 410 74 590 90
rect 410 54 449 74
rect 74 40 168 54
rect -130 24 168 40
rect 196 49 304 54
rect 332 49 449 54
rect 196 40 449 49
rect 483 40 517 74
rect 551 54 590 74
rect 551 40 630 54
rect 196 24 630 40
<< polycont >>
rect 237 182 271 212
rect 237 104 271 134
rect -74 40 -40 74
rect 40 40 74 74
rect 449 40 483 74
rect 517 40 551 74
<< corelocali >>
rect 144 301 168 331
rect 196 301 356 331
rect 144 255 356 273
rect 144 254 304 255
rect -86 211 -17 245
rect 17 227 86 245
rect 17 211 35 227
rect -86 193 35 211
rect 69 193 86 227
rect 144 220 168 254
rect 196 245 304 254
rect 196 237 208 245
tri 208 237 216 245 nw
tri 201 230 208 237 nw
rect 300 221 304 245
rect 332 221 356 255
rect 144 219 190 220
tri 190 219 191 220 nw
rect 300 219 356 221
rect 414 227 586 245
tri 223 212 228 217 se
rect 228 212 272 217
tri 212 201 223 212 se
rect 223 201 237 212
rect -86 177 86 193
tri 202 191 212 201 se
rect 212 191 237 201
rect -86 143 -17 177
rect 17 155 86 177
rect 116 175 144 191
tri 193 182 202 191 se
rect 202 182 237 191
rect 271 182 272 212
rect 17 143 35 155
rect -86 121 35 143
rect 69 121 86 155
tri 185 174 193 182 se
rect 193 175 272 182
rect 193 174 225 175
tri 225 174 226 175 nw
tri 172 161 185 174 se
rect 185 161 212 174
tri 212 161 225 174 nw
rect 116 125 144 141
rect -86 107 86 121
rect 172 97 200 161
tri 200 149 212 161 nw
tri 290 149 300 159 se
rect 300 149 328 219
rect 414 193 431 227
rect 465 226 586 227
rect 465 193 483 226
rect 414 192 483 193
rect 517 192 586 226
rect 356 175 384 191
tri 283 142 290 149 se
rect 290 147 328 149
rect 290 142 323 147
tri 323 142 328 147 nw
tri 282 141 283 142 se
rect 283 141 322 142
tri 322 141 323 142 nw
rect 414 158 586 192
rect 414 155 483 158
rect 232 134 305 141
rect 232 104 237 134
rect 271 124 305 134
tri 305 124 322 141 nw
rect 356 125 384 141
rect 271 119 300 124
tri 300 119 305 124 nw
rect 414 121 431 155
rect 465 124 483 155
rect 517 124 586 158
rect 465 121 586 124
rect 271 104 280 119
rect 232 99 280 104
tri 280 99 300 119 nw
rect 414 107 586 121
rect 144 96 200 97
rect -90 40 -74 74
rect -40 66 40 74
rect -40 40 -17 66
rect 17 40 40 66
rect 74 40 90 74
rect 144 62 168 96
tri 316 95 318 97 se
rect 318 95 356 97
rect 196 71 200 79
tri 292 71 304 83 se
rect 196 62 304 71
rect 144 61 304 62
rect 332 61 356 95
rect 144 43 356 61
rect 433 74 567 77
rect 433 40 449 74
rect 551 40 567 74
rect 433 37 567 40
rect 144 -15 168 15
rect 196 -15 356 15
<< viali >>
rect 35 193 69 227
rect 35 121 69 155
rect 113 174 147 175
rect 113 142 116 174
rect 116 142 144 174
rect 144 142 147 174
rect 113 141 147 142
rect 431 193 465 227
rect 353 174 387 175
rect 353 142 356 174
rect 356 142 384 174
rect 384 142 387 174
rect 353 141 387 142
rect 431 121 465 155
rect -17 32 17 66
rect 483 40 517 74
<< metal1 >>
rect 28 227 76 316
rect 116 263 144 316
rect 190 287 238 345
rect 28 207 35 227
rect 0 193 35 207
rect 69 207 76 227
rect 104 207 144 263
rect 69 193 144 207
rect 0 185 144 193
rect 0 179 156 185
rect 0 159 104 179
rect 28 155 76 159
rect 28 121 35 155
rect 69 121 76 155
rect 104 126 156 127
tri 104 121 109 126 ne
rect 109 121 156 126
rect 28 116 76 121
tri 28 90 54 116 ne
rect 54 102 76 116
tri 76 102 88 114 sw
tri -23 78 -19 82 se
rect -19 78 19 82
tri 19 78 23 82 sw
tri -26 75 -23 78 se
rect -23 75 23 78
tri 23 75 26 78 sw
rect -26 21 26 23
tri -26 20 -25 21 ne
rect -25 20 25 21
tri 25 20 26 21 nw
tri -25 14 -19 20 ne
rect -19 14 19 20
tri 19 14 25 20 nw
rect 54 0 88 102
rect 116 -15 144 121
rect 200 0 228 287
rect 272 29 300 316
rect 356 263 384 316
rect 344 257 396 263
rect 424 227 472 316
rect 424 207 431 227
rect 396 205 431 207
rect 344 198 431 205
rect 347 193 431 198
rect 465 207 472 227
rect 465 193 500 207
rect 347 175 500 193
rect 347 141 353 175
rect 387 159 500 175
rect 387 141 393 159
rect 347 129 393 141
tri 347 127 349 129 ne
rect 349 127 391 129
tri 391 127 393 129 nw
rect 424 155 472 159
rect 262 -29 310 29
rect 356 -15 384 127
rect 424 121 431 155
rect 465 122 472 155
rect 465 121 470 122
rect 424 120 470 121
tri 470 120 472 122 nw
tri 412 108 424 120 se
rect 424 108 458 120
tri 458 108 470 120 nw
rect 412 0 446 108
tri 446 96 458 108 nw
tri 474 84 478 88 se
rect 478 84 522 88
tri 522 84 526 88 sw
rect 474 82 526 84
rect 474 20 526 30
tri 474 14 480 20 ne
rect 480 14 520 20
tri 520 14 526 20 nw
<< via1 >>
rect 104 175 156 179
rect 104 141 113 175
rect 113 141 147 175
rect 147 141 156 175
rect 104 127 156 141
rect -26 66 26 75
rect -26 32 -17 66
rect -17 32 17 66
rect 17 32 26 66
rect -26 23 26 32
rect 344 205 396 257
rect 474 74 526 82
rect 474 40 483 74
rect 483 40 517 74
rect 517 40 526 74
rect 474 30 526 40
<< metal2 >>
rect -130 213 344 257
rect 321 205 344 213
rect 396 205 630 257
rect -130 127 104 179
rect 156 171 188 179
rect 156 127 630 171
rect -130 82 630 93
rect -130 75 474 82
rect -130 59 -26 75
rect -32 24 -26 59
rect 26 59 474 75
rect 26 24 32 59
rect 526 59 630 82
rect 474 24 526 30
<< labels >>
flabel metal1 s 272 208 300 244 0 FreeSans 100 90 0 0 br
flabel metal1 s 200 208 228 244 0 FreeSans 100 0 0 0 bl
flabel metal2 s 592 217 623 251 0 FreeSans 2000 0 0 0 vdd
flabel metal2 s -122 138 -91 172 0 FreeSans 2000 0 0 0 gnd
flabel metal2 s 234 59 265 93 0 FreeSans 2000 0 0 0 wl
flabel nbase s 358 31 368 41 0 FreeSans 40 90 0 0 VPB
port 1 nsew
flabel pwell s 132 34 142 46 0 FreeSans 100 90 0 0 VNB
port 0 nsew
<< properties >>
string GDS_FILE sky130_fd_bd_sram__openram_cell_6t_dummy.gds
string GDS_END 13168
string GDS_START 170
string path -2.250 1.425 2.250 1.425 
<< end >>
