VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colend_met2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colend_met2 ;
  ORIGIN 0.055 -0.020 ;
  SIZE 1.310 BY 2.035 ;
  OBS
      LAYER met1 ;
        RECT 1.070 1.695 1.255 1.955 ;
        RECT -0.055 0.745 0.130 1.005 ;
      LAYER met2 ;
        RECT 0.000 1.955 1.200 2.055 ;
        RECT 0.000 1.695 1.255 1.955 ;
        RECT 0.000 1.600 1.200 1.695 ;
        RECT 0.000 1.180 1.200 1.460 ;
        RECT 0.000 1.005 1.200 1.030 ;
        RECT -0.055 0.745 1.200 1.005 ;
        RECT 0.000 0.580 1.200 0.745 ;
        RECT 0.000 0.020 1.200 0.405 ;
  END
END sky130_fd_bd_sram__sram_sp_colend_met2
END LIBRARY

