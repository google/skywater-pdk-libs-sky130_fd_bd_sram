VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_cell
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_cell ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.200 BY 1.580 ;
  OBS
      LAYER nwell ;
        RECT 0.720 0.000 1.200 1.580 ;
      LAYER li1 ;
        RECT 0.190 1.505 0.330 1.580 ;
        RECT 0.535 0.910 0.705 1.060 ;
        RECT 0.000 0.710 0.070 0.870 ;
        RECT 1.115 0.705 1.200 0.875 ;
        RECT 0.535 0.520 0.705 0.670 ;
        RECT 0.190 0.000 0.330 0.075 ;
      LAYER met1 ;
        RECT 1.115 0.705 1.200 0.875 ;
  END
END sky130_fd_bd_sram__openram_sp_cell
END LIBRARY

