# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_blkinv_opt2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_blkinv_opt2 ;
  ORIGIN  0.055000  0.505000 ;
  SIZE  3.165000 BY  1.475000 ;
  OBS
    LAYER li1 ;
      RECT 0.090000 -0.125000 0.260000  0.775000 ;
      RECT 0.510000 -0.015000 1.300000  0.155000 ;
      RECT 0.510000  0.155000 0.680000  0.790000 ;
      RECT 0.860000  0.335000 2.405000  0.480000 ;
      RECT 0.860000  0.480000 2.155000  0.530000 ;
      RECT 0.860000  0.530000 1.650000  0.585000 ;
      RECT 0.860000  0.585000 1.110000  0.665000 ;
      RECT 1.080000 -0.415000 1.250000 -0.245000 ;
      RECT 1.480000  0.260000 2.155000  0.310000 ;
      RECT 1.480000  0.310000 2.405000  0.335000 ;
      RECT 2.295000  0.000000 2.635000  0.050000 ;
      RECT 2.295000  0.050000 2.880000  0.170000 ;
      RECT 2.295000  0.620000 2.880000  0.740000 ;
      RECT 2.295000  0.740000 2.635000  0.790000 ;
      RECT 2.495000  0.170000 2.880000  0.190000 ;
      RECT 2.495000  0.600000 2.880000  0.620000 ;
      RECT 2.585000  0.190000 2.880000  0.265000 ;
      RECT 2.585000  0.265000 3.055000  0.525000 ;
      RECT 2.585000  0.525000 2.880000  0.600000 ;
    LAYER mcon ;
      RECT 1.980000 0.310000 2.150000 0.480000 ;
      RECT 2.465000 0.000000 2.635000 0.085000 ;
      RECT 2.465000 0.705000 2.635000 0.790000 ;
      RECT 2.970000 0.310000 3.055000 0.480000 ;
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000  0.000000 ;
      RECT -0.055000  0.000000 0.390000  0.130000 ;
      RECT -0.055000  0.660000 0.390000  0.790000 ;
      RECT -0.055000  0.790000 0.130000  0.845000 ;
      RECT  0.000000  0.130000 0.390000  0.660000 ;
      RECT  0.590000  0.000000 0.840000  0.790000 ;
      RECT  1.035000 -0.505000 1.295000 -0.155000 ;
      RECT  1.040000  0.000000 1.290000  0.790000 ;
      RECT  1.490000  0.000000 1.740000  0.790000 ;
      RECT  1.935000  0.220000 2.195000  0.570000 ;
      RECT  1.940000  0.000000 2.190000  0.220000 ;
      RECT  1.940000  0.570000 2.190000  0.790000 ;
      RECT  2.435000  0.000000 3.110000  0.130000 ;
      RECT  2.435000  0.130000 3.055000  0.660000 ;
      RECT  2.435000  0.660000 3.110000  0.790000 ;
      RECT  2.925000 -0.055000 3.110000  0.000000 ;
      RECT  2.925000  0.790000 3.110000  0.845000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 -0.040000 ;
      RECT -0.055000 -0.040000 0.140000  0.000000 ;
      RECT -0.055000  0.000000 0.240000  0.130000 ;
      RECT -0.055000  0.660000 0.240000  0.790000 ;
      RECT -0.055000  0.790000 0.140000  0.830000 ;
      RECT -0.055000  0.830000 0.130000  0.845000 ;
      RECT -0.040000  0.130000 0.240000  0.140000 ;
      RECT -0.040000  0.650000 0.240000  0.660000 ;
      RECT  0.000000  0.140000 0.240000  0.650000 ;
      RECT  1.600000  0.000000 3.110000  0.130000 ;
      RECT  1.600000  0.130000 3.055000  0.660000 ;
      RECT  1.600000  0.660000 3.110000  0.790000 ;
      RECT  2.925000 -0.055000 3.110000  0.000000 ;
      RECT  2.925000  0.790000 3.110000  0.845000 ;
    LAYER met3 ;
      RECT -0.040000 -0.040000 0.140000 0.000000 ;
      RECT -0.040000  0.000000 3.055000 0.140000 ;
      RECT -0.040000  0.650000 3.055000 0.790000 ;
      RECT -0.040000  0.790000 0.140000 0.830000 ;
      RECT  0.000000  0.140000 3.055000 0.205000 ;
      RECT  0.000000  0.205000 0.205000 0.585000 ;
      RECT  0.000000  0.585000 3.055000 0.650000 ;
    LAYER nwell ;
      RECT 0.000000 0.000000 1.755000 0.790000 ;
      RECT 0.320000 0.790000 1.610000 0.970000 ;
    LAYER via ;
      RECT 2.925000 0.660000 3.110000 0.845000 ;
    LAYER via2 ;
      RECT -0.040000 -0.040000 0.140000 0.140000 ;
  END
END sky130_fd_bd_sram__sram_dp_blkinv_opt2
END LIBRARY
