# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_colend_swldrv_opt1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_colend_swldrv_opt1 ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  3.165000 BY  1.980000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1.310000 0.085000 ;
      RECT 0.000000 0.085000 1.180000 0.385000 ;
      RECT 0.000000 0.385000 0.165000 0.545000 ;
      RECT 0.000000 0.975000 3.055000 1.145000 ;
      RECT 2.295000 0.585000 3.055000 0.975000 ;
      RECT 2.300000 0.000000 2.635000 0.085000 ;
      RECT 2.300000 0.310000 2.470000 0.480000 ;
      RECT 2.835000 0.120000 3.005000 0.270000 ;
    LAYER mcon ;
      RECT 0.000000 0.200000 0.085000 0.370000 ;
      RECT 2.465000 0.000000 2.635000 0.085000 ;
      RECT 2.970000 0.775000 3.055000 0.945000 ;
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.185000 0.130000 ;
      RECT -0.055000  1.565000 0.185000 1.825000 ;
      RECT  0.000000  0.130000 0.185000 1.565000 ;
      RECT  0.000000  1.825000 0.185000 1.925000 ;
      RECT  0.590000  0.000000 0.840000 1.925000 ;
      RECT  1.040000  0.000000 1.290000 1.925000 ;
      RECT  1.490000  0.000000 1.740000 1.925000 ;
      RECT  1.940000  0.000000 2.190000 1.925000 ;
      RECT  2.435000  0.000000 3.110000 0.130000 ;
      RECT  2.435000  0.130000 3.055000 0.730000 ;
      RECT  2.435000  0.730000 3.110000 0.990000 ;
      RECT  2.435000  0.990000 3.055000 1.925000 ;
      RECT  2.925000 -0.055000 3.110000 0.000000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 -0.040000 ;
      RECT -0.055000 -0.040000 0.140000  0.000000 ;
      RECT -0.055000  0.000000 0.240000  0.130000 ;
      RECT -0.055000  1.565000 3.055000  1.825000 ;
      RECT -0.040000  0.130000 0.240000  0.140000 ;
      RECT  0.000000  0.140000 0.240000  0.240000 ;
      RECT  0.000000  1.470000 3.055000  1.565000 ;
      RECT  0.000000  1.825000 3.055000  1.925000 ;
      RECT  1.600000  0.000000 3.110000  0.130000 ;
      RECT  1.600000  0.130000 3.055000  0.730000 ;
      RECT  1.600000  0.730000 3.110000  0.990000 ;
      RECT  1.600000  0.990000 3.055000  1.085000 ;
      RECT  2.925000 -0.055000 3.110000  0.000000 ;
    LAYER met3 ;
      RECT -0.040000 -0.040000 0.140000 0.000000 ;
      RECT -0.040000  0.000000 3.055000 0.140000 ;
      RECT  0.000000  0.140000 3.055000 0.205000 ;
    LAYER nwell ;
      RECT 0.000000 0.375000 1.755000 0.785000 ;
    LAYER nwell ;
      RECT 1.510000 0.160000 1.755000 0.375000 ;
    LAYER nwell ;
      RECT 1.575000 0.000000 1.755000 0.160000 ;
    LAYER pwell ;
      RECT 0.000000 0.000000 1.575000 0.160000 ;
    LAYER pwell ;
      RECT 0.000000 0.160000 1.510000 0.375000 ;
    LAYER pwell ;
      RECT 0.000000 0.915000 3.055000 1.205000 ;
    LAYER pwell ;
      RECT 2.095000 0.000000 2.595000 0.715000 ;
      RECT 2.095000 0.715000 3.055000 0.915000 ;
    LAYER via ;
      RECT 2.925000 0.730000 3.110000 0.990000 ;
    LAYER via2 ;
      RECT -0.040000 -0.040000 0.140000 0.140000 ;
  END
END sky130_fd_bd_sram__sram_dp_colend_swldrv_opt1
END LIBRARY
