magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1202 -1320 2236 1738
<< nwell >>
rect 412 -60 976 478
<< pwell >>
rect 58 100 142 136
<< nmos >>
rect 196 266 344 296
rect 196 194 344 224
<< pmos >>
rect 582 272 806 302
rect 582 182 806 212
<< ndiff >>
rect 196 348 344 369
rect 196 314 257 348
rect 291 314 344 348
rect 196 296 344 314
rect 196 224 344 266
rect 196 176 344 194
rect 196 142 259 176
rect 293 142 344 176
rect 196 134 344 142
<< pdiff >>
rect 582 348 806 369
rect 582 314 677 348
rect 711 314 806 348
rect 582 302 806 314
rect 582 260 806 272
rect 582 226 677 260
rect 711 226 806 260
rect 582 212 806 226
rect 582 170 806 182
rect 582 136 677 170
rect 711 136 806 170
rect 582 128 806 136
<< ndiffc >>
rect 257 314 291 348
rect 259 142 293 176
<< pdiffc >>
rect 677 314 711 348
rect 677 226 711 260
rect 677 136 711 170
<< psubdiff >>
rect 58 135 142 136
rect 58 101 83 135
rect 117 101 142 135
rect 58 100 142 101
<< nsubdiff >>
rect 861 171 899 196
rect 861 137 863 171
rect 897 137 899 171
rect 861 112 899 137
<< psubdiffcont >>
rect 83 101 117 135
<< nsubdiffcont >>
rect 863 137 897 171
<< poly >>
rect 76 316 130 332
rect 76 282 86 316
rect 120 296 130 316
rect 460 296 582 302
rect 120 282 196 296
rect 76 266 196 282
rect 344 272 582 296
rect 806 272 832 302
rect 344 266 478 272
rect 76 208 196 224
rect 76 174 86 208
rect 120 194 196 208
rect 344 212 490 224
rect 344 194 582 212
rect 120 174 130 194
rect 76 158 130 174
rect 458 182 582 194
rect 806 182 832 212
<< polycont >>
rect 86 282 120 316
rect 86 174 120 208
<< locali >>
rect 70 282 86 316
rect 120 282 136 316
rect 210 314 257 348
rect 291 314 677 348
rect 711 314 888 348
rect 70 174 86 208
rect 120 174 136 208
rect 208 142 254 176
rect 293 142 340 176
rect 509 170 543 314
rect 660 226 677 260
rect 711 226 727 260
rect 845 171 915 172
rect 509 169 598 170
rect 660 169 677 170
rect 509 136 677 169
rect 711 136 728 170
rect 845 137 863 171
rect 897 137 915 171
rect 845 136 915 137
rect 66 135 142 136
rect 66 101 83 135
rect 117 101 142 135
rect 509 135 685 136
rect 509 134 572 135
rect 66 100 142 101
<< viali >>
rect 254 142 259 176
rect 259 142 288 176
rect 677 226 711 260
rect 863 137 897 171
rect 83 101 117 135
<< metal1 >>
rect 246 176 294 402
rect 76 136 124 148
rect 246 142 254 176
rect 288 142 294 176
rect 246 136 294 142
rect 76 135 294 136
rect 76 101 83 135
rect 117 101 294 135
rect 76 100 294 101
rect 76 88 124 100
rect 246 29 294 100
rect 670 260 720 402
rect 670 226 677 260
rect 711 226 720 260
rect 670 170 720 226
rect 845 171 912 178
rect 845 170 863 171
rect 670 137 863 170
rect 897 137 912 171
rect 670 136 912 137
rect 670 30 720 136
rect 849 128 912 136
<< labels >>
rlabel corelocali s 103 191 103 191 4 B
rlabel corelocali s 103 299 103 299 4 A
rlabel corelocali s 854 331 854 331 4 Z
rlabel metal1 s 696 94 696 94 4 VDD
port 1 nsew
rlabel metal1 s 268 82 268 82 4 GND
port 0 nsew
<< properties >>
string FIXED_BBOX 58 53 915 396
string GDS_FILE sky130_fd_bd_sram__openram_nand2_dec.gds
string GDS_END 4008
string GDS_START 162
<< end >>
