magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1260 1500 1418
<< pdiff >>
rect 38 118 80 158
rect 38 0 80 40
<< viali >>
rect 0 62 17 96
<< metal1 >>
rect 0 117 42 158
rect 0 0 42 41
<< via1 >>
rect -11 96 26 105
rect -11 62 0 96
rect 0 62 17 96
rect 17 62 26 96
rect -11 53 26 62
use sky130_fd_bd_sram__sram_dp_horstrap_half  sky130_fd_bd_sram__sram_dp_horstrap_half_0
timestamp 0
transform 1 0 0 0 1 0
box 0 0 240 158
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_horstrap_half1.gds
string GDS_END 2296
string GDS_START 1908
<< end >>
