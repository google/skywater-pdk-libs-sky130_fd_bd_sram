* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_cell_6t VNB VPB VPB
X0 VPB a_146_104# a_146_182# VPB sky130_fd_pr__pfet_01v8_hvt w=140000u l=150000u
X1 a_146_182# wl a_146_182# VPB sky130_fd_pr__pfet_01v8_hvt w=70000u l=95000u
X2 bl wl a_146_104# SUBS sky130_fd_pr__special_nfet_latch w=140000u l=150000u
X3 gnd a_146_104# a_146_182# SUBS sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X4 a_146_104# a_146_182# gnd SUBS sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X5 a_146_104# wl a_146_104# VPB sky130_fd_pr__pfet_01v8_hvt w=70000u l=95000u
X6 a_146_182# wl br SUBS sky130_fd_pr__special_nfet_latch w=140000u l=150000u
X7 a_146_104# a_146_182# VPB VPB sky130_fd_pr__pfet_01v8_hvt w=140000u l=150000u
.ends
