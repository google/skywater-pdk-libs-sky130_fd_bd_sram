VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_corner_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_corner_ce ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.300 BY 2.055 ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 0.445 2.055 ;
      LAYER li1 ;
        RECT 0.000 1.160 1.300 1.875 ;
        RECT 0.000 0.990 0.340 1.160 ;
        RECT 0.520 0.810 1.130 0.990 ;
        RECT 0.000 0.275 1.130 0.810 ;
        RECT 0.160 0.000 1.130 0.275 ;
      LAYER mcon ;
        RECT 0.285 1.610 0.455 1.780 ;
        RECT 0.285 1.250 0.455 1.420 ;
        RECT 0.790 0.755 0.960 0.925 ;
        RECT 0.900 0.055 1.070 0.225 ;
      LAYER met1 ;
        RECT 0.000 1.025 0.090 2.055 ;
        RECT 0.250 1.205 0.550 2.055 ;
        POLYGON 0.250 1.205 0.310 1.205 0.310 1.145 ;
        POLYGON 0.090 1.105 0.170 1.025 0.090 1.025 ;
        RECT 0.000 0.730 0.170 1.025 ;
        RECT 0.000 0.000 0.070 0.730 ;
        POLYGON 0.070 0.730 0.170 0.730 0.070 0.630 ;
        POLYGON 0.310 0.495 0.310 0.395 0.210 0.395 ;
        RECT 0.310 0.395 0.550 1.205 ;
        RECT 0.210 0.170 0.550 0.395 ;
        RECT 0.210 0.000 0.380 0.170 ;
        POLYGON 0.380 0.170 0.550 0.170 0.380 0.000 ;
        RECT 0.760 1.215 1.060 2.055 ;
        RECT 0.760 0.365 0.990 1.215 ;
        POLYGON 0.990 1.215 1.060 1.215 0.990 1.145 ;
        POLYGON 0.990 0.465 1.090 0.365 0.990 0.365 ;
        RECT 0.760 0.160 1.090 0.365 ;
        POLYGON 0.760 0.160 0.865 0.160 0.865 0.055 ;
        RECT 0.865 0.055 1.090 0.160 ;
        POLYGON 0.865 0.055 0.920 0.055 0.920 0.000 ;
        RECT 0.920 0.000 1.090 0.055 ;
  END
END sky130_fd_bd_sram__sram_sp_corner_ce
END LIBRARY

