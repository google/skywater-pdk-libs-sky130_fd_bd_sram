* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_dp_nand4_dec A B C D GND VDD Z
X0 a_406_159# C a_406_87# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 Z A VDD VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 VDD D a_1166_91# VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_406_231# B a_406_159# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_406_303# B VDD VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 VDD C a_406_303# VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 a_406_303# A a_406_231# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_406_87# D GND GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
