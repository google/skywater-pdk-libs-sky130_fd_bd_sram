magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1260 1751 1418
<< pdiff >>
rect 38 118 80 158
rect 400 118 442 158
rect 38 0 80 40
rect 400 0 442 40
use sky130_fd_bd_sram__sram_dp_horstrap_half2  sky130_fd_bd_sram__sram_dp_horstrap_half2_0
timestamp 0
transform 1 0 0 0 1 0
box -11 0 240 158
use sky130_fd_bd_sram__sram_dp_horstrap_p1m_siz  sky130_fd_bd_sram__sram_dp_horstrap_p1m_siz_0
timestamp 0
transform 1 0 0 0 1 0
box 0 24 480 135
use sky130_fd_bd_sram__sram_dp_horstrap_npsdm  sky130_fd_bd_sram__sram_dp_horstrap_npsdm_0
timestamp 0
transform 1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_horstrap_limcon  sky130_fd_bd_sram__sram_dp_horstrap_limcon_0
timestamp 0
transform 1 0 0 0 -1 158
box 14 0 466 158
use sky130_fd_bd_sram__sram_dp_horstrap_half1  sky130_fd_bd_sram__sram_dp_horstrap_half1_0
timestamp 0
transform -1 0 480 0 1 0
box -11 0 240 158
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_horstrap2a.gds
string GDS_END 6354
string GDS_START 5930
<< end >>
