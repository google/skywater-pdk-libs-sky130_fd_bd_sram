VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_rowend_replica
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_rowend_replica ;
  ORIGIN 0.055 0.000 ;
  SIZE 1.355 BY 1.580 ;
  PIN VPWR
    ANTENNADIFFAREA 0.021600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.705 0.085 0.875 ;
      LAYER met1 ;
        RECT 0.000 1.315 0.070 1.580 ;
        RECT 0.000 1.285 0.130 1.315 ;
        RECT -0.055 1.025 0.130 1.285 ;
        RECT 0.000 0.990 0.130 1.025 ;
        RECT 0.000 0.635 0.105 0.990 ;
        RECT 0.000 0.000 0.070 0.635 ;
      LAYER met2 ;
        RECT -0.055 1.025 1.300 1.285 ;
    END
  END VPWR
  PIN WL
    PORT
      LAYER li1 ;
        RECT 0.395 0.200 0.905 0.370 ;
      LAYER mcon ;
        RECT 0.565 0.200 0.735 0.370 ;
      LAYER met1 ;
        POLYGON 0.540 0.440 0.540 0.420 0.520 0.420 ;
        RECT 0.540 0.420 0.760 0.440 ;
        POLYGON 0.760 0.440 0.780 0.420 0.760 0.420 ;
        RECT 0.520 0.100 0.780 0.420 ;
        POLYGON 0.520 0.100 0.550 0.100 0.550 0.070 ;
        RECT 0.550 0.070 0.750 0.100 ;
        POLYGON 0.750 0.100 0.780 0.100 0.750 0.070 ;
      LAYER via ;
        RECT 0.520 0.150 0.780 0.410 ;
      LAYER met2 ;
        RECT 0.000 0.295 1.300 0.465 ;
        RECT 0.520 0.120 0.780 0.295 ;
    END
  END WL
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 1.300 1.580 ;
      LAYER li1 ;
        RECT 0.305 0.965 0.475 1.135 ;
        RECT 0.565 0.960 0.735 1.130 ;
        RECT 0.305 0.605 0.475 0.775 ;
        RECT 0.565 0.620 0.735 0.790 ;
      LAYER met1 ;
        RECT 0.270 0.610 0.510 1.580 ;
        RECT 0.270 0.600 0.500 0.610 ;
        POLYGON 0.500 0.610 0.510 0.610 0.500 0.600 ;
        RECT 0.790 0.610 1.030 1.580 ;
        POLYGON 0.790 0.610 0.800 0.610 0.800 0.600 ;
        RECT 0.800 0.600 1.030 0.610 ;
        POLYGON 0.270 0.600 0.270 0.540 0.210 0.540 ;
        RECT 0.270 0.540 0.380 0.600 ;
        RECT 0.210 0.000 0.380 0.540 ;
        POLYGON 0.380 0.600 0.500 0.600 0.380 0.480 ;
        POLYGON 0.800 0.600 0.920 0.600 0.920 0.480 ;
        RECT 0.920 0.540 1.030 0.600 ;
        POLYGON 1.030 0.600 1.090 0.540 1.030 0.540 ;
        RECT 0.920 0.000 1.090 0.540 ;
      LAYER met2 ;
        RECT 0.000 0.635 1.300 0.855 ;
  END
END sky130_fd_bd_sram__openram_sp_rowend_replica
END LIBRARY

