# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_cell_met23_opt1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_cell_met23_opt1 ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  2.510000 BY  1.580000 ;
  OBS
    LAYER met1 ;
      RECT -0.055000 0.660000 0.130000 0.920000 ;
      RECT  2.270000 0.660000 2.455000 0.920000 ;
    LAYER met2 ;
      RECT -0.055000 0.660000 2.455000 0.920000 ;
      RECT  0.000000 0.120000 2.400000 0.360000 ;
      RECT  0.000000 0.600000 2.400000 0.660000 ;
      RECT  0.000000 0.920000 2.400000 0.980000 ;
      RECT  0.000000 1.220000 2.400000 1.460000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 2.400000 0.205000 ;
      RECT 0.000000 0.505000 2.400000 1.075000 ;
      RECT 0.000000 1.375000 2.400000 1.580000 ;
  END
END sky130_fd_bd_sram__sram_dp_cell_met23_opt1
END LIBRARY
