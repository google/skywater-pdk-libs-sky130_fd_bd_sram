
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.SUBCKT sky130_fd_bd_sram__openram_cell_6t bl br wl vdd gnd
* Inverter 1
Xsky130_fd_pr__special_nfet_latch_bar Qbar Q gnd gnd sky130_fd_pr__special_nfet_latch W=0.210 L=0.150
Xsky130_fd_pr__special_pfet_latch_bar Qbar Q vdd vdd sky130_fd_pr__special_pfet_latch W=0.140 L=0.150

* Inverer 2
Xsky130_fd_pr__special_nfet_latch_tru Q Qbar gnd gnd sky130_fd_pr__special_nfet_latch W=0.210 L=0.150 
Xsky130_fd_pr__special_pfet_latch_tru Q Qbar vdd vdd sky130_fd_pr__special_pfet_latch W=0.140 L=0.150

* Access transistors
Xspecial_nfet_pass_tru bl wl Q gnd special_nfet_pass W=0.140 L=0.150
Xspecial_nfet_pass_bar br wl Qbar gnd special_nfet_pass W=0.140 L=0.150

* Parasitic transistors
Xpdo_tru Q wl Q vdd sky130_fd_pr__special_pfet_latch W=0.140 L=0.025
Xpdo_bar Qbar wl Qbar vdd sky130_fd_pr__special_pfet_latch W=0.140 L=0.025

.ENDS sky130_fd_bd_sram__openram_cell_6t
