magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1246 -1260 1455 1309
use sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos  sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos_0
timestamp 0
transform 1 0 14 0 1 0
box 0 0 1 1
use sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos  sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos_1
timestamp 0
transform 1 0 14 0 1 48
box 0 0 1 1
use sky130_fd_bd_sram__openram_sp_cell_fom_serif_pmos  sky130_fd_bd_sram__openram_sp_cell_fom_serif_pmos_0
timestamp 0
transform 1 0 194 0 1 48
box 0 0 1 1
use sky130_fd_bd_sram__openram_sp_cell_fom_serif_pmos  sky130_fd_bd_sram__openram_sp_cell_fom_serif_pmos_1
timestamp 0
transform 1 0 194 0 1 0
box 0 0 1 1
<< properties >>
string GDS_FILE sky130_fd_bd_sram__openram_sp_cell_fom_serifs.gds
string GDS_END 782
string GDS_START 482
<< end >>
