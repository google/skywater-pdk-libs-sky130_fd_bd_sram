* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


* Top level circuit sky130_fd_bd_sram__openram_cell_1rw_1r_dummy
X0 a_38_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X1 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X2 a_400_n79# gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch w=105000u l=185000u
X3 br0 wl0 a_400_291# gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X4 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch w=105000u l=185000u
X5 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch w=105000u l=185000u
X6 gnd gnd a_400_133# gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X7 a_400_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X8 a_38_n79# gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch w=105000u l=185000u
X9 bl0 wl0 a_38_291# gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X10 a_400_133# wl1 br1 gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X11 gnd gnd a_38_133# gnd sky130_fd_pr__special_nfet_latch w=210000u l=150000u
.end
