* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




.subckt sky130_fd_bd_sram__sram_sp_cell_opt1 bl br vgnd vnb vpb vpwr wl
Xsky130_fd_bd_sram__sram_sp_cell_opt1_ce_0 vgnd bl a_70_79# vnb vpwr a_62_220# wl
+ vpb br a_108_24# sky130_fd_bd_sram__sram_sp_cell_opt1_ce
.ends
