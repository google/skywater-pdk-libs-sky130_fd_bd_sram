# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell_metopt1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell_metopt1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.200000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.705000 0.085000 0.875000 ;
      RECT 0.335000 1.495000 0.505000 1.580000 ;
      RECT 0.695000 0.000000 0.865000 0.085000 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
    LAYER met1 ;
      POLYGON 1.085000 0.645000 1.095000 0.645000 1.095000 0.635000 ;
      RECT 0.000000 0.000000 0.070000 0.605000 ;
      RECT 0.000000 0.605000 0.130000 0.925000 ;
      RECT 0.000000 0.925000 0.070000 1.580000 ;
      RECT 0.300000 1.435000 0.540000 1.580000 ;
      RECT 0.350000 0.000000 0.490000 1.435000 ;
      RECT 0.660000 0.000000 0.900000 0.145000 ;
      RECT 0.710000 0.145000 0.850000 1.580000 ;
      RECT 1.070000 0.990000 1.200000 1.315000 ;
      RECT 1.085000 0.645000 1.200000 0.990000 ;
      RECT 1.095000 0.635000 1.200000 0.645000 ;
      RECT 1.130000 0.000000 1.200000 0.635000 ;
      RECT 1.130000 1.315000 1.200000 1.580000 ;
  END
END sky130_fd_bd_sram__sram_sp_cell_metopt1
END LIBRARY
