magic
tech sky130A
magscale 1 2
timestamp 1621288235
<< dnwell >>
rect 0 0 260 411
<< pwell >>
rect -26 80 286 362
<< psubdiff >>
rect 0 201 260 336
rect 0 167 79 201
rect 113 167 147 201
rect 181 167 260 201
rect 0 142 260 167
rect 17 108 243 142
rect 0 106 260 108
<< psubdiffcont >>
rect 79 167 113 201
rect 147 167 181 201
rect 0 108 17 142
rect 243 108 260 142
<< poly >>
rect 0 24 260 54
<< locali >>
rect 0 341 70 375
rect 104 341 260 375
rect 0 303 260 341
rect 0 269 70 303
rect 104 269 260 303
rect 0 235 260 269
rect 0 167 79 201
rect 113 167 147 201
rect 181 167 260 201
rect 0 162 260 167
rect 0 142 158 162
rect 17 128 158 142
rect 192 142 260 162
rect 192 128 243 142
rect 17 108 243 128
rect 0 90 260 108
rect 0 56 158 90
rect 192 56 260 90
rect 0 55 260 56
rect 27 3 240 55
<< viali >>
rect 70 341 104 375
rect 70 269 104 303
rect 158 128 192 162
rect 158 56 192 90
<< metal1 >>
rect 0 337 30 411
rect 0 204 18 337
tri 18 325 30 337 nw
rect 62 375 110 411
rect 62 341 70 375
rect 104 341 110 375
tri 50 311 62 323 se
rect 62 311 110 341
rect 50 303 110 311
rect 50 269 70 303
rect 104 269 110 303
rect 50 231 110 269
tri 18 204 34 220 sw
tri 50 219 62 231 ne
rect 0 146 34 204
rect 0 0 14 146
tri 14 126 34 146 nw
tri 42 76 62 96 se
rect 62 76 110 231
rect 42 34 110 76
rect 42 0 76 34
tri 76 0 110 34 nw
rect 150 311 198 411
rect 230 337 260 411
tri 230 325 242 337 ne
tri 198 311 210 323 sw
rect 150 231 210 311
rect 150 162 198 231
tri 198 219 210 231 nw
rect 150 128 158 162
rect 192 128 198 162
rect 150 90 198 128
tri 226 205 242 221 se
rect 242 205 260 337
rect 226 146 260 205
tri 226 126 246 146 ne
rect 150 56 158 90
rect 192 76 198 90
tri 198 76 218 96 sw
rect 192 56 218 76
rect 150 34 218 56
tri 150 0 184 34 ne
rect 184 0 218 34
rect 246 0 260 146
<< end >>
