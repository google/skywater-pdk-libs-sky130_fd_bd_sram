VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_cell_metopt1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_cell_metopt1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.200 BY 1.580 ;
  OBS
      LAYER li1 ;
        RECT 0.335 1.495 0.505 1.580 ;
        RECT 0.000 0.705 0.085 0.875 ;
        RECT 1.115 0.705 1.200 0.875 ;
        RECT 0.695 0.000 0.865 0.085 ;
      LAYER met1 ;
        RECT 0.000 0.925 0.070 1.580 ;
        RECT 0.300 1.435 0.540 1.580 ;
        RECT 0.000 0.605 0.130 0.925 ;
        RECT 0.000 0.000 0.070 0.605 ;
        RECT 0.350 0.000 0.490 1.435 ;
        RECT 0.710 0.145 0.850 1.580 ;
        RECT 1.130 1.315 1.200 1.580 ;
        RECT 1.070 0.990 1.200 1.315 ;
        RECT 1.085 0.645 1.200 0.990 ;
        POLYGON 1.085 0.645 1.095 0.645 1.095 0.635 ;
        RECT 1.095 0.635 1.200 0.645 ;
        RECT 0.660 0.000 0.900 0.145 ;
        RECT 1.130 0.000 1.200 0.635 ;
  END
END sky130_fd_bd_sram__openram_sp_cell_metopt1
END LIBRARY

