VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colenda_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colenda_ce ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.200 BY 2.055 ;
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 0.480 2.055 ;
      LAYER pwell ;
        RECT 0.700 0.530 1.200 1.680 ;
      LAYER li1 ;
        RECT 0.000 1.175 1.200 1.875 ;
        RECT 0.000 0.990 0.340 1.175 ;
        RECT 0.520 0.810 1.200 1.005 ;
        RECT 0.000 0.275 1.200 0.810 ;
        RECT 0.335 0.075 0.505 0.085 ;
        RECT 0.070 0.000 1.130 0.075 ;
      LAYER mcon ;
        RECT 0.335 0.000 0.505 0.085 ;
      LAYER met1 ;
        RECT 0.000 1.025 0.090 2.055 ;
        RECT 0.305 1.590 0.485 2.055 ;
        POLYGON 0.305 1.590 0.345 1.590 0.345 1.550 ;
        POLYGON 0.090 1.105 0.170 1.025 0.090 1.025 ;
        RECT 0.000 0.730 0.170 1.025 ;
        RECT 0.000 0.000 0.070 0.730 ;
        POLYGON 0.070 0.730 0.170 0.730 0.070 0.630 ;
        RECT 0.345 0.145 0.485 1.590 ;
        RECT 0.710 1.595 0.890 2.055 ;
        RECT 0.300 0.000 0.540 0.145 ;
        RECT 0.710 0.000 0.850 1.595 ;
        POLYGON 0.850 1.595 0.890 1.595 0.850 1.555 ;
        RECT 1.050 1.595 1.200 2.055 ;
        POLYGON 1.050 1.595 1.090 1.595 1.090 1.555 ;
        RECT 1.090 1.555 1.200 1.595 ;
        POLYGON 1.090 1.555 1.130 1.555 1.130 1.515 ;
        RECT 1.130 0.000 1.200 1.555 ;
  END
END sky130_fd_bd_sram__sram_sp_colenda_ce
END LIBRARY

