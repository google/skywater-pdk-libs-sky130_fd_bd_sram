# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_cell
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_cell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.710000 0.085000 0.870000 ;
      RECT 0.210000 0.000000 0.380000 0.085000 ;
      RECT 0.210000 0.310000 0.380000 0.480000 ;
      RECT 0.210000 1.100000 0.380000 1.270000 ;
      RECT 0.210000 1.495000 0.380000 1.580000 ;
      RECT 0.535000 0.910000 0.695000 0.940000 ;
      RECT 0.545000 0.770000 0.695000 0.910000 ;
      RECT 0.875000 0.725000 1.010000 0.895000 ;
      RECT 1.280000 0.300000 1.420000 0.470000 ;
      RECT 1.280000 0.705000 1.420000 0.875000 ;
      RECT 1.280000 1.110000 1.420000 1.280000 ;
      RECT 1.705000 0.640000 1.865000 0.670000 ;
      RECT 1.705000 0.670000 1.855000 0.810000 ;
      RECT 2.020000 0.000000 2.190000 0.085000 ;
      RECT 2.020000 0.310000 2.190000 0.480000 ;
      RECT 2.020000 1.100000 2.190000 1.270000 ;
      RECT 2.020000 1.495000 2.190000 1.580000 ;
      RECT 2.315000 0.710000 2.400000 0.870000 ;
    LAYER nwell ;
      RECT 0.720000 0.000000 1.680000 1.580000 ;
  END
END sky130_fd_bd_sram__sram_dp_cell
END LIBRARY
