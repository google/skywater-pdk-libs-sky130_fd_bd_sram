magic
tech sky130A
magscale 1 2
timestamp 1621288248
<< dnwell >>
rect 0 0 260 316
<< nwell >>
rect 0 0 260 316
<< pdiff >>
rect 14 142 27 174
rect 233 142 246 174
<< pdiffc >>
rect 0 142 14 174
rect 246 142 260 174
<< nsubdiff >>
rect 83 226 177 252
rect 83 192 113 226
rect 147 192 177 226
rect 83 158 177 192
rect 83 124 113 158
rect 147 124 177 158
rect 83 100 177 124
<< nsubdiffcont >>
rect 113 192 147 226
rect 113 124 147 158
<< poly >>
rect 0 262 260 292
rect 40 90 73 262
rect 187 90 220 262
rect 40 74 220 90
rect 40 54 79 74
rect 0 40 79 54
rect 113 40 147 74
rect 181 54 220 74
rect 181 40 260 54
rect 0 24 260 40
<< polycont >>
rect 79 40 113 74
rect 147 40 181 74
<< corelocali >>
rect 44 227 216 245
rect 44 193 61 227
rect 95 226 216 227
rect 95 193 113 226
rect 44 192 113 193
rect 147 192 216 226
rect 0 175 14 191
rect 44 158 216 192
rect 246 175 260 191
rect 44 155 113 158
rect 0 125 14 141
rect 44 121 61 155
rect 95 124 113 155
rect 147 124 216 158
rect 246 125 260 141
rect 95 121 216 124
rect 44 107 216 121
rect 63 74 197 77
rect 63 40 79 74
rect 181 40 197 74
rect 63 37 197 40
<< viali >>
rect 61 193 95 227
rect 0 174 17 175
rect 0 142 14 174
rect 14 142 17 174
rect 0 141 17 142
rect 61 121 95 155
rect 243 174 260 175
rect 243 142 246 174
rect 246 142 260 174
rect 243 141 260 142
rect 113 40 147 74
<< metal1 >>
rect 0 263 14 316
rect 0 256 26 263
rect 25 206 26 256
rect 0 198 26 206
rect 54 227 102 316
rect 0 175 23 198
rect 17 141 23 175
rect 0 129 23 141
rect 0 127 21 129
tri 21 127 23 129 nw
rect 54 193 61 227
rect 95 193 102 227
rect 54 155 102 193
rect 0 0 14 127
rect 54 121 61 155
rect 95 122 102 155
rect 95 121 100 122
rect 54 120 100 121
tri 100 120 102 122 nw
rect 158 122 206 316
rect 246 263 260 316
rect 234 256 260 263
rect 234 206 235 256
rect 234 198 260 206
rect 237 175 260 198
rect 237 141 243 175
rect 237 129 260 141
tri 237 127 239 129 ne
rect 239 127 260 129
tri 42 108 54 120 se
rect 54 108 76 120
rect 42 0 76 108
tri 76 96 100 120 nw
tri 158 96 184 122 ne
rect 184 108 206 122
tri 206 108 218 120 sw
tri 104 84 108 88 se
rect 108 84 152 88
tri 152 84 156 88 sw
rect 104 81 156 84
rect 104 31 105 81
rect 155 31 156 81
rect 104 20 156 31
tri 104 14 110 20 ne
rect 110 14 150 20
tri 150 14 156 20 nw
rect 184 0 218 108
rect 246 0 260 127
<< via1 >>
rect -10 206 25 256
rect 235 206 270 256
rect 105 74 155 81
rect 105 40 113 74
rect 113 40 147 74
rect 147 40 155 74
rect 105 31 155 40
<< end >>
