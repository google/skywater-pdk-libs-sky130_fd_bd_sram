# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell_via
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell_via ;
  ORIGIN  0.055000 -0.635000 ;
  SIZE  1.310000 BY  0.650000 ;
  OBS
    LAYER met1 ;
      RECT -0.055000 0.635000 0.130000 0.895000 ;
      RECT  1.070000 1.025000 1.255000 1.285000 ;
    LAYER met2 ;
      RECT -0.055000 0.635000 0.130000 0.895000 ;
      RECT  1.070000 1.025000 1.255000 1.285000 ;
  END
END sky130_fd_bd_sram__sram_sp_cell_via
END LIBRARY
