* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* SPICE3 file created from sky130_fd_bd_sram__openram_dff.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_dff D Q CLK VDD GND
M1000 a_511_725# a_n8_115# VDD VDD pshort W=3 L=0.15 m=1 mult=1
M1001 a_353_115# CLK a_11_624# GND nshort W=1 L=0.15 m=1 mult=1
M1002 a_353_725# a_203_89# a_11_624# VDD pshort W=3 L=0.15 m=1 mult=1
M1003 a_11_624# a_203_89# a_161_115# GND nshort W=1 L=0.15 m=1 mult=1
M1004 a_11_624# CLK a_161_725# VDD pshort W=3 L=0.15 m=1 mult=1
M1005 GND Q a_703_115# GND nshort W=1 L=0.15 m=1 mult=1
M1006 VDD Q a_703_725# VDD pshort W=3 L=0.15 m=1 mult=1
M1007 a_203_89# CLK GND GND nshort W=1 L=0.15 m=1 mult=1
M1008 a_203_89# CLK VDD VDD pshort W=3 L=0.15 m=1 mult=1
M1009 a_161_115# D GND GND nshort W=1 L=0.15 m=1 mult=1
M1010 a_161_725# D VDD VDD pshort W=3 L=0.15 m=1 mult=1
M1011 GND a_11_624# a_n8_115# GND nshort W=1 L=0.15 m=1 mult=1
M1012 a_703_115# a_203_89# ON GND nshort W=1 L=0.15 m=1 mult=1
M1013 VDD a_11_624# a_n8_115# VDD pshort W=3 L=0.15 m=1 mult=1
M1014 a_703_725# CLK ON VDD pshort W=3 L=0.15 m=1 mult=1
M1015 Q ON VDD VDD pshort W=3 L=0.15 m=1 mult=1
M1016 Q ON GND GND nshort W=1 L=0.15 m=1 mult=1
M1017 ON a_203_89# a_511_725# VDD pshort W=3 L=0.15 m=1 mult=1
M1018 ON CLK a_511_115# GND nshort W=1 L=0.15 m=1 mult=1
M1019 GND a_n8_115# a_353_115# GND nshort W=1 L=0.15 m=1 mult=1
M1020 VDD a_n8_115# a_353_725# VDD pshort W=3 L=0.15 m=1 mult=1
M1021 a_511_115# a_n8_115# GND GND nshort W=1 L=0.15 m=1 mult=1
.ends
