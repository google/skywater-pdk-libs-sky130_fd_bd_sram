magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1330 -1320 2582 1734
<< nwell >>
rect 414 -60 1322 474
<< pwell >>
rect -64 260 -10 343
<< nmos >>
rect 128 250 276 280
rect 128 178 276 208
rect 128 106 276 136
<< pmos >>
rect 584 206 808 236
rect 584 106 808 136
rect 1016 106 1240 136
<< ndiff >>
rect 128 327 276 351
rect 128 293 191 327
rect 225 293 276 327
rect 128 280 276 293
rect 128 208 276 250
rect 128 136 276 178
rect 128 95 276 106
rect 128 61 189 95
rect 223 61 276 95
rect 128 53 276 61
<< pdiff >>
rect 584 288 808 296
rect 584 254 679 288
rect 713 254 808 288
rect 584 236 808 254
rect 584 188 808 206
rect 584 154 679 188
rect 713 154 808 188
rect 584 136 808 154
rect 1016 188 1240 204
rect 1016 154 1111 188
rect 1145 154 1240 188
rect 1016 136 1240 154
rect 584 95 808 106
rect 584 61 679 95
rect 713 61 808 95
rect 584 46 808 61
rect 1016 95 1240 106
rect 1016 61 1111 95
rect 1145 61 1240 95
rect 1016 46 1240 61
<< ndiffc >>
rect 191 293 225 327
rect 189 61 223 95
<< pdiffc >>
rect 679 254 713 288
rect 679 154 713 188
rect 1111 154 1145 188
rect 679 61 713 95
rect 1111 61 1145 95
<< psubdiff >>
rect -64 318 -10 343
rect -64 284 -54 318
rect -20 284 -10 318
rect -64 260 -10 284
<< nsubdiff >>
rect 1086 288 1110 322
rect 1144 288 1170 322
<< psubdiffcont >>
rect -54 284 -20 318
<< nsubdiffcont >>
rect 1110 288 1144 322
<< poly >>
rect 46 300 100 316
rect 46 266 56 300
rect 90 280 100 300
rect 331 300 386 316
rect 331 280 342 300
rect 90 266 128 280
rect 46 250 128 266
rect 276 266 342 280
rect 376 266 386 300
rect 928 300 982 316
rect 276 250 386 266
rect -64 210 -10 226
rect -64 176 -54 210
rect -20 208 -10 210
rect 928 266 938 300
rect 972 266 982 300
rect 470 208 584 236
rect -20 178 128 208
rect 276 206 584 208
rect 808 206 834 236
rect 928 234 982 266
rect 276 178 500 206
rect -20 176 -10 178
rect -64 160 -10 176
rect 940 136 970 234
rect 46 120 128 136
rect 46 86 56 120
rect 90 106 128 120
rect 276 106 584 136
rect 808 106 834 136
rect 940 106 1016 136
rect 1240 106 1266 136
rect 90 86 100 106
rect 46 70 100 86
<< polycont >>
rect 56 266 90 300
rect 342 266 376 300
rect -54 176 -20 210
rect 938 266 972 300
rect 56 86 90 120
<< locali >>
rect -54 334 180 368
rect -54 318 -20 334
rect 140 330 180 334
rect 140 327 272 330
rect -54 260 -20 284
rect 40 266 56 300
rect 90 266 106 300
rect 140 293 184 327
rect 225 293 272 327
rect 1110 322 1148 338
rect 140 291 272 293
rect 326 300 411 302
rect 326 255 342 300
rect 376 260 411 300
rect 922 300 1007 302
rect 511 288 687 289
rect 376 255 394 260
rect 326 243 394 255
rect 511 255 679 288
rect -70 176 -54 210
rect -20 176 -4 210
rect 40 86 56 120
rect 90 86 106 120
rect 511 95 545 255
rect 662 254 679 255
rect 713 254 730 288
rect 922 255 938 300
rect 972 260 1007 300
rect 1145 288 1148 322
rect 1110 272 1148 288
rect 972 255 990 260
rect 922 243 990 255
rect 662 154 679 188
rect 713 154 1111 188
rect 1145 154 1161 188
rect 142 61 189 95
rect 223 61 679 95
rect 713 61 1111 95
rect 1145 61 1322 95
<< viali >>
rect 184 293 191 327
rect 191 293 218 327
rect 342 266 376 289
rect 342 255 376 266
rect 938 266 972 289
rect 938 255 972 266
rect 1111 288 1144 322
rect 1144 288 1145 322
rect 679 154 713 188
rect 1111 154 1145 188
<< metal1 >>
rect 178 327 224 368
rect 178 293 184 327
rect 218 293 224 327
rect 178 -44 224 293
rect 326 290 394 302
rect 326 289 395 290
rect 326 286 342 289
rect 376 286 395 289
rect 326 234 334 286
rect 386 234 395 286
rect 326 227 395 234
rect 672 188 720 368
rect 1104 322 1152 368
rect 922 290 990 302
rect 922 289 991 290
rect 922 286 938 289
rect 972 286 991 289
rect 922 234 930 286
rect 982 234 991 286
rect 922 227 991 234
rect 1104 288 1111 322
rect 1145 288 1152 322
rect 672 154 679 188
rect 713 154 720 188
rect 672 14 720 154
rect 1104 188 1152 288
rect 1104 154 1111 188
rect 1145 154 1152 188
rect 1104 14 1152 154
<< via1 >>
rect 334 255 342 286
rect 342 255 376 286
rect 376 255 386 286
rect 334 234 386 255
rect 930 255 938 286
rect 938 255 972 286
rect 972 255 982 286
rect 930 234 982 255
<< metal2 >>
rect 326 286 1009 288
rect 326 234 334 286
rect 386 260 930 286
rect 386 234 395 260
rect 326 227 395 234
rect 922 234 930 260
rect 982 260 1009 286
rect 982 234 991 260
rect 922 227 991 234
<< labels >>
rlabel metal1 s 677 338 715 356 4 VDD
port 1 nsew
rlabel metal1 s 1109 338 1147 356 4 VDD
port 1 nsew
rlabel corelocali s 1294 78 1294 78 4 Z
rlabel corelocali s 70 284 70 284 4 C
rlabel metal1 s 183 338 219 356 4 GND
port 0 nsew
rlabel corelocali s -40 196 -40 196 4 B
rlabel corelocali s 70 106 70 106 4 A
<< properties >>
string FIXED_BBOX -72 35 1321 351
string GDS_FILE sky130_fd_bd_sram__openram_nand3_dec.gds
string GDS_END 6070
string GDS_START 162
<< end >>
