# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_opt4bi
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_opt4bi ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  3.165000 BY  1.690000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.165000 1.300000 0.270000 ;
      RECT 0.000000 0.270000 0.650000 0.435000 ;
      RECT 0.000000 1.170000 0.315000 1.580000 ;
      RECT 0.510000 0.000000 0.680000 0.055000 ;
      RECT 0.510000 0.055000 1.300000 0.165000 ;
      RECT 0.510000 1.175000 1.435000 1.490000 ;
      RECT 0.540000 0.685000 2.790000 0.895000 ;
      RECT 0.540000 0.895000 1.495000 0.950000 ;
      RECT 1.480000 0.185000 2.155000 0.505000 ;
      RECT 2.295000 0.000000 2.635000 0.160000 ;
      RECT 2.295000 0.160000 2.490000 0.535000 ;
      RECT 2.295000 1.045000 2.490000 1.420000 ;
      RECT 2.295000 1.420000 2.635000 1.580000 ;
      RECT 2.630000 0.320000 2.985000 0.465000 ;
      RECT 2.630000 0.465000 2.790000 0.685000 ;
      RECT 2.630000 0.895000 2.790000 1.115000 ;
      RECT 2.630000 1.115000 2.985000 1.260000 ;
      RECT 2.780000 0.090000 2.985000 0.120000 ;
      RECT 2.780000 0.120000 3.005000 0.270000 ;
      RECT 2.780000 0.270000 2.985000 0.320000 ;
      RECT 2.780000 1.260000 2.985000 1.490000 ;
      RECT 2.930000 0.625000 3.055000 0.955000 ;
    LAYER mcon ;
      RECT 0.050000 1.255000 0.220000 1.425000 ;
      RECT 0.175000 0.215000 0.345000 0.385000 ;
      RECT 0.630000 1.270000 0.800000 1.440000 ;
      RECT 1.530000 0.260000 1.700000 0.430000 ;
      RECT 2.465000 0.000000 2.635000 0.085000 ;
      RECT 2.465000 1.495000 2.635000 1.580000 ;
      RECT 2.490000 0.705000 2.660000 0.875000 ;
      RECT 2.970000 0.705000 3.055000 0.875000 ;
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.390000 0.130000 ;
      RECT  0.000000  0.130000 0.390000 0.475000 ;
      RECT  0.000000  0.475000 0.185000 0.680000 ;
      RECT  0.000000  1.140000 0.370000 1.580000 ;
      RECT  0.585000  1.180000 0.845000 1.530000 ;
      RECT  0.590000  0.000000 0.840000 1.180000 ;
      RECT  0.590000  1.530000 0.840000 1.580000 ;
      RECT  1.040000  0.000000 1.290000 1.580000 ;
      RECT  1.485000  0.170000 1.745000 0.520000 ;
      RECT  1.490000  0.000000 1.740000 0.170000 ;
      RECT  1.490000  0.520000 1.740000 1.580000 ;
      RECT  1.940000  0.000000 2.190000 1.580000 ;
      RECT  2.370000  0.600000 2.790000 1.020000 ;
      RECT  2.375000  0.535000 2.790000 0.600000 ;
      RECT  2.435000  0.000000 3.110000 0.130000 ;
      RECT  2.435000  0.130000 3.055000 0.355000 ;
      RECT  2.435000  1.200000 3.055000 1.450000 ;
      RECT  2.435000  1.450000 3.110000 1.580000 ;
      RECT  2.925000 -0.055000 3.110000 0.000000 ;
      RECT  2.925000  1.580000 3.110000 1.635000 ;
      RECT  2.970000  0.355000 3.055000 1.200000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 -0.040000 ;
      RECT -0.055000 -0.040000 0.140000  0.000000 ;
      RECT -0.055000  0.000000 0.240000  0.130000 ;
      RECT -0.040000  0.130000 0.240000  0.140000 ;
      RECT  0.000000  0.140000 0.240000  0.240000 ;
      RECT  0.000000  0.480000 2.080000  0.905000 ;
      RECT  0.025000  1.145000 0.345000  1.580000 ;
      RECT  1.600000  0.000000 3.110000  0.130000 ;
      RECT  1.600000  0.130000 3.055000  0.185000 ;
      RECT  1.600000  0.185000 2.080000  0.480000 ;
      RECT  1.600000  0.905000 2.080000  1.395000 ;
      RECT  1.600000  1.395000 3.055000  1.450000 ;
      RECT  1.600000  1.450000 3.110000  1.580000 ;
      RECT  2.370000  0.605000 3.055000  0.845000 ;
      RECT  2.370000  0.845000 2.780000  0.925000 ;
      RECT  2.925000 -0.055000 3.110000  0.000000 ;
      RECT  2.925000  1.580000 3.110000  1.635000 ;
    LAYER met3 ;
      RECT -0.040000 -0.040000 0.140000 0.000000 ;
      RECT -0.040000  0.000000 3.055000 0.140000 ;
      RECT  0.000000  0.140000 3.055000 0.205000 ;
      RECT  0.000000  0.505000 3.055000 1.075000 ;
      RECT  0.000000  1.375000 3.055000 1.580000 ;
    LAYER nwell ;
      RECT 0.000000 0.000000 1.755000 1.580000 ;
    LAYER pwell ;
      RECT 2.095000 1.380000 2.595000 1.580000 ;
    LAYER via ;
      RECT 0.055000 1.220000 0.315000 1.480000 ;
      RECT 2.445000 0.635000 2.705000 0.895000 ;
      RECT 2.925000 1.450000 3.110000 1.635000 ;
    LAYER via2 ;
      RECT -0.040000 -0.040000 0.140000 0.140000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_opt4bi
END LIBRARY
