# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.200000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      POLYGON 0.305000 1.150000 0.355000 1.150000 0.305000 1.100000 ;
      POLYGON 0.930000 0.475000 0.930000 0.415000 0.870000 0.415000 ;
      RECT 0.000000 0.710000 0.070000 0.870000 ;
      RECT 0.190000 0.000000 0.330000 0.075000 ;
      RECT 0.190000 0.310000 0.330000 0.395000 ;
      RECT 0.190000 0.395000 0.350000 0.480000 ;
      RECT 0.190000 1.100000 0.305000 1.150000 ;
      RECT 0.190000 1.150000 0.355000 1.185000 ;
      RECT 0.190000 1.185000 0.330000 1.270000 ;
      RECT 0.190000 1.505000 0.330000 1.580000 ;
      RECT 0.535000 0.520000 0.705000 0.670000 ;
      RECT 0.535000 0.910000 0.705000 1.060000 ;
      RECT 0.870000 0.305000 1.010000 0.415000 ;
      RECT 0.870000 1.105000 1.010000 1.275000 ;
      RECT 0.930000 0.415000 1.010000 0.475000 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
    LAYER met1 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
    LAYER nwell ;
      RECT 0.690000 0.065000 1.200000 1.515000 ;
      RECT 0.720000 0.000000 1.200000 0.065000 ;
      RECT 0.720000 1.515000 1.200000 1.580000 ;
  END
END sky130_fd_bd_sram__sram_sp_cell
END LIBRARY
