magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1302 -1315 1884 1631
<< poly >>
rect 410 341 624 371
rect 410 103 624 133
rect 428 25 624 55
rect 428 -25 478 25
rect 428 -55 624 -25
<< metal2 >>
rect -42 323 624 371
rect 438 309 520 323
rect -42 261 404 275
rect 554 261 624 275
rect -42 213 624 261
rect -42 199 404 213
rect 554 199 624 213
rect 438 151 520 165
rect -42 103 624 151
rect -42 -55 624 55
<< labels >>
flabel metal2 s 225 222 256 256 0 FreeSans 2000 0 0 0 gnd
flabel metal2 s 224 -14 255 19 0 FreeSans 2000 0 0 0 gnd
flabel metal2 s 324 331 355 365 0 FreeSans 2000 0 0 0 wl0
flabel metal2 s 303 107 335 141 0 FreeSans 2000 0 0 0 wl1
<< properties >>
string FIXED_BBOX 0 0 624 395
string GDS_FILE sky130_fd_bd_sram__openram_cell_1rw_1r_cap_row.gds
string GDS_END 4434
string GDS_START 182
<< end >>
