# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_horstrap_limcon
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_horstrap_limcon ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  2.260000 BY  0.790000 ;
  OBS
    LAYER li1 ;
      RECT 0.070000 0.000000 1.670000 0.075000 ;
      RECT 0.070000 0.665000 0.590000 0.790000 ;
      RECT 0.490000 0.075000 1.670000 0.125000 ;
      RECT 0.730000 0.665000 1.910000 0.715000 ;
      RECT 0.730000 0.715000 2.330000 0.790000 ;
      RECT 1.810000 0.000000 2.330000 0.125000 ;
    LAYER mcon ;
      RECT 0.395000 0.705000 0.565000 0.790000 ;
      RECT 0.755000 0.705000 0.925000 0.790000 ;
      RECT 1.475000 0.000000 1.645000 0.085000 ;
      RECT 1.835000 0.000000 2.005000 0.085000 ;
    LAYER met1 ;
      RECT 0.395000 0.705000 0.565000 0.790000 ;
      RECT 0.755000 0.705000 0.925000 0.790000 ;
      RECT 1.475000 0.000000 1.645000 0.085000 ;
      RECT 1.835000 0.000000 2.005000 0.085000 ;
  END
END sky130_fd_bd_sram__sram_dp_horstrap_limcon
END LIBRARY
