
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.SUBCKT sky130_fd_bd_sram__openram_cell_1rw_1r bl0 br0 bl1 br1 wl0 wl1 vdd gnd
** N=11 EP=8 IP=0 FDC=16
*.SEEDPROM

* Bitcell Core
X0 Q wl1 bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X1 gnd Q_bar Q gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X2 gnd Q_bar Q gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X3 bl0 wl0 Q gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X4 Q_bar wl1 br1 gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X5 gnd Q Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X6 gnd Q Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X7 br0 wl0 Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.15u m=1
X8 vdd Q Q_bar vdd sky130_fd_pr__special_pfet_latch W=0.14u L=0.15u m=1
X9 Q Q_bar vdd vdd sky130_fd_pr__special_pfet_latch W=0.14u L=0.15u m=1

* drainOnly PMOS
X10 Q_bar wl1 Q_bar vdd sky130_fd_pr__special_pfet_latch W=0.14u L=0.08u m=1
X11 Q wl0 Q vdd sky130_fd_pr__special_pfet_latch W=0.14u L=0.08u m=1

* drainOnly NMOS
X12 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.08u m=1
X14 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch W=0.21u L=0.08u m=1

.ENDS
