magic
tech sky130A
magscale 1 2
timestamp 1623356714
<< nwell >>
rect 594 -79 1502 437
<< pwell >>
rect 115 289 223 343
<< nmos >>
rect 308 229 456 259
rect 308 157 456 187
rect 308 85 456 115
<< pmos >>
rect 764 185 988 215
rect 764 85 988 115
rect 1196 85 1420 115
<< ndiff >>
rect 308 333 456 342
rect 308 299 364 333
rect 405 299 456 333
rect 308 259 456 299
rect 308 187 456 229
rect 308 115 456 157
rect 308 74 456 85
rect 308 40 369 74
rect 403 40 456 74
rect 308 32 456 40
<< pdiff >>
rect 764 267 988 275
rect 764 233 859 267
rect 893 233 988 267
rect 764 215 988 233
rect 764 167 988 185
rect 764 133 859 167
rect 893 133 988 167
rect 764 115 988 133
rect 1196 167 1420 183
rect 1196 133 1291 167
rect 1325 133 1420 167
rect 1196 115 1420 133
rect 764 74 988 85
rect 764 40 859 74
rect 893 40 988 74
rect 764 27 988 40
rect 1196 74 1420 85
rect 1196 40 1291 74
rect 1325 40 1420 74
rect 1196 28 1420 40
<< ndiffc >>
rect 364 299 405 333
rect 369 40 403 74
<< pdiffc >>
rect 859 233 893 267
rect 859 133 893 167
rect 1291 133 1325 167
rect 859 40 893 74
rect 1291 40 1325 74
<< psubdiff >>
rect 115 333 223 343
rect 115 299 139 333
rect 173 299 223 333
rect 115 289 223 299
<< nsubdiff >>
rect 1266 237 1290 271
rect 1324 237 1350 271
<< psubdiffcont >>
rect 139 299 173 333
<< nsubdiffcont >>
rect 1290 237 1324 271
<< poly >>
rect 511 279 566 295
rect 511 259 522 279
rect 6 243 308 259
rect 6 209 16 243
rect 50 229 308 243
rect 456 245 522 259
rect 556 245 566 279
rect 1108 279 1162 295
rect 456 229 566 245
rect 50 209 61 229
rect 6 193 61 209
rect 1108 245 1118 279
rect 1152 245 1162 279
rect 650 187 764 215
rect 116 171 308 187
rect 116 137 126 171
rect 160 157 308 171
rect 456 185 764 187
rect 988 185 1014 215
rect 1108 213 1162 245
rect 456 157 680 185
rect 160 137 170 157
rect 116 121 170 137
rect 1120 115 1150 213
rect 226 99 308 115
rect 226 65 236 99
rect 270 85 308 99
rect 456 85 764 115
rect 988 85 1014 115
rect 1120 85 1196 115
rect 1420 85 1446 115
rect 270 65 280 85
rect 226 49 280 65
<< polycont >>
rect 16 209 50 243
rect 522 245 556 279
rect 1118 245 1152 279
rect 126 137 160 171
rect 236 65 270 99
<< locali >>
rect 115 299 139 333
rect 173 299 364 333
rect 405 299 453 333
rect 506 279 591 281
rect 0 209 16 243
rect 50 209 66 243
rect 506 234 522 279
rect 556 239 591 279
rect 1102 279 1187 281
rect 691 267 867 268
rect 556 234 574 239
rect 506 222 574 234
rect 691 234 859 267
rect 110 137 126 171
rect 160 137 176 171
rect 220 65 236 99
rect 270 65 286 99
rect 691 74 725 234
rect 842 233 859 234
rect 893 233 910 267
rect 1102 234 1118 279
rect 1152 239 1187 279
rect 1290 271 1328 287
rect 1152 234 1170 239
rect 1102 222 1170 234
rect 1324 237 1328 271
rect 1290 204 1328 237
rect 842 133 859 167
rect 893 133 1291 167
rect 1325 133 1341 167
rect 322 40 369 74
rect 403 40 859 74
rect 893 40 1291 74
rect 1325 40 1502 74
<< viali >>
rect 364 299 398 333
rect 522 245 556 268
rect 522 234 556 245
rect 1118 245 1152 268
rect 1118 234 1152 245
rect 1290 237 1324 271
rect 859 133 893 167
rect 1291 133 1325 167
<< metal1 >>
rect 358 333 404 349
rect 358 299 364 333
rect 398 299 404 333
rect 358 -63 404 299
rect 506 269 574 281
rect 506 268 575 269
rect 506 265 522 268
rect 556 265 575 268
rect 506 213 514 265
rect 566 213 575 265
rect 506 206 575 213
rect 852 167 900 347
rect 1102 269 1170 281
rect 1284 271 1332 302
rect 1102 268 1171 269
rect 1102 265 1118 268
rect 1152 265 1171 268
rect 1102 213 1110 265
rect 1162 213 1171 265
rect 1102 206 1171 213
rect 1284 237 1290 271
rect 1324 237 1332 271
rect 852 133 859 167
rect 893 133 900 167
rect 852 -7 900 133
rect 1284 167 1332 237
rect 1284 133 1291 167
rect 1325 133 1332 167
rect 1284 -7 1332 133
<< via1 >>
rect 514 234 522 265
rect 522 234 556 265
rect 556 234 566 265
rect 514 213 566 234
rect 1110 234 1118 265
rect 1118 234 1152 265
rect 1152 234 1162 265
rect 1110 213 1162 234
<< metal2 >>
rect 506 265 575 267
rect 506 213 514 265
rect 566 213 575 265
rect 506 211 575 213
rect 1102 265 1189 267
rect 1102 213 1110 265
rect 1162 239 1189 265
rect 1162 213 1171 239
rect 1102 211 1171 213
rect 506 159 1171 211
<< labels >>
rlabel metal1 s 358 -63 404 349 4 GND
rlabel locali s 1474 57 1474 57 4 Z
rlabel metal1 s 381 141 381 141 4 gnd
rlabel metal1 s 852 -7 900 347 4 VDD
rlabel metal1 s 1284 -7 1332 302 4 VDD
rlabel metal1 s 876 170 876 170 4 vdd
rlabel metal1 s 1308 147 1308 147 4 vdd
rlabel metal1 s 381 143 381 143 4 gnd
rlabel polycont 253 82 253 82 1 A
rlabel polycont 143 154 143 154 1 B
rlabel polycont 33 226 33 226 1 C
<< properties >>
string FIXED_BBOX 0 0 1502 316
<< end >>
