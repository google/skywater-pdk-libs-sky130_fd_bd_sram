# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_cell_1rw_1r_cap_col
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_cell_1rw_1r_cap_col ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.120000 BY  2.370000 ;
  OBS
    LAYER met1 ;
      RECT 0.390000 0.000000 0.570000 2.370000 ;
      RECT 0.750000 0.000000 0.930000 2.370000 ;
      RECT 1.070000 0.790000 1.330000 1.500000 ;
      RECT 1.110000 0.000000 1.290000 0.790000 ;
      RECT 1.110000 1.500000 1.290000 2.370000 ;
      RECT 1.470000 0.000000 1.650000 2.370000 ;
      RECT 1.830000 0.000000 2.010000 2.370000 ;
    LAYER met2 ;
      RECT 0.000000 0.870000 3.120000 1.420000 ;
    LAYER via ;
      RECT 1.070000 1.020000 1.330000 1.280000 ;
  END
END sky130_fd_bd_sram__openram_cell_1rw_1r_cap_col
END LIBRARY
