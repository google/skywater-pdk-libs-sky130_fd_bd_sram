magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1256 -1260 1265 1261
use sky130_fd_bd_sram__sram_dp_cell_poly_srf_opta  sky130_fd_bd_sram__sram_dp_cell_poly_srf_opta_0
timestamp 0
transform -1 0 5 0 1 0
box 0 0 1 1
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_wls_p1m_ser.gds
string GDS_END 532
string GDS_START 312
<< end >>
