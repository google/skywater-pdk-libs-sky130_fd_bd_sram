# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.005000 BY  0.005000 ;
END sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta
END LIBRARY
