VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_cell_addpoly
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_cell_addpoly ;
  ORIGIN 0.000 -0.120 ;
  SIZE 0.080 BY 1.340 ;
END sky130_fd_bd_sram__openram_sp_cell_addpoly
END LIBRARY

