# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_rowendb
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_rowendb ;
  ORIGIN  0.000000  0.055000 ;
  SIZE  1.115000 BY  1.635000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 0.415000 1.580000 ;
      RECT 0.775000 0.000000 0.940000 0.545000 ;
      RECT 0.775000 1.170000 0.940000 1.580000 ;
    LAYER mcon ;
      RECT 0.050000 0.000000 0.220000 0.085000 ;
      RECT 0.855000 0.200000 0.940000 0.370000 ;
    LAYER met1 ;
      RECT 0.005000  0.000000 0.265000 0.130000 ;
      RECT 0.045000  0.130000 0.225000 1.580000 ;
      RECT 0.445000  0.000000 0.995000 0.130000 ;
      RECT 0.445000  0.130000 0.940000 0.680000 ;
      RECT 0.445000  0.680000 1.115000 0.940000 ;
      RECT 0.445000  0.940000 0.730000 1.580000 ;
      RECT 0.810000 -0.055000 0.995000 0.000000 ;
    LAYER met2 ;
      RECT 0.445000  0.000000 0.995000  0.130000 ;
      RECT 0.445000  0.130000 0.980000  0.140000 ;
      RECT 0.445000  0.140000 0.940000  0.240000 ;
      RECT 0.800000 -0.040000 0.995000  0.000000 ;
      RECT 0.810000 -0.055000 0.995000 -0.040000 ;
    LAYER met3 ;
      RECT 0.445000  0.000000 0.980000 0.140000 ;
      RECT 0.445000  0.140000 0.940000 0.205000 ;
      RECT 0.445000  1.375000 0.940000 1.580000 ;
      RECT 0.800000 -0.040000 0.980000 0.000000 ;
    LAYER nwell ;
      RECT 0.605000 0.000000 0.940000 1.580000 ;
    LAYER pwell ;
      RECT 0.185000 0.000000 0.475000 1.580000 ;
    LAYER via2 ;
      RECT 0.800000 -0.040000 0.980000 0.140000 ;
  END
END sky130_fd_bd_sram__sram_dp_rowendb
END LIBRARY
