
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* SPICE3 file created from sky130_fd_bd_sram__openram_sram_dff.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_sram_dff D Q clk vdd gnd
X1000 a_511_725# a_n8_115# vdd vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1001 a_353_115# clk a_11_624# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1002 a_353_725# a_203_89# a_11_624# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1003 a_11_624# a_203_89# a_161_115# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1004 a_11_624# clk a_161_725# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1005 gnd Q a_703_115# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1006 vdd Q a_703_725# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1007 a_203_89# clk gnd gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1008 a_203_89# clk vdd vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1009 a_161_115# D gnd gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1010 a_161_725# D vdd vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1011 gnd a_11_624# a_n8_115# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1012 a_703_115# a_203_89# ON gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1013 vdd a_11_624# a_n8_115# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1014 a_703_725# clk ON vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1015 Q ON vdd vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1016 Q ON gnd gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1017 ON a_203_89# a_511_725# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1018 ON clk a_511_115# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1019 gnd a_n8_115# a_353_115# gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
X1020 vdd a_n8_115# a_353_725# vdd sky130_fd_pr__pfet_01v8 W=3u L=0.15u m=1
X1021 a_511_115# a_n8_115# gnd gnd sky130_fd_pr__nfet_01v8 W=1u L=0.15u m=1
.ends
