magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE sky130_fd_bd_sram__openram_sp_cell_fom_serif_pmos.gds
string GDS_END 258
string GDS_START 190
<< end >>
