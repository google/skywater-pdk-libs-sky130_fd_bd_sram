* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_sense_amp" ******************************

.SUBCKT sky130_fd_bd_sram__openram_sense_amp BL BR DOUT EN VDD GND
M1000 GND EN a_56_432# GND nshort W=0.65 L=0.15 m=1 mult=1
M1001 a_56_432# dint_bar dint GND nshort W=0.65 L=0.15 m=1 mult=1
M1002 dint_bar dint a_56_432# GND nshort W=0.65 L=0.15 m=1 mult=1

M1003 VDD dint_bar dint VDD pshort W=1.26 L=0.15 m=1 mult=1
M1004 dint_bar dint VDD VDD pshort W=1.26 L=0.15 m=1 mult=1

M1005 BL EN dint VDD pshort W=2 L=0.15 m=1 mult=1
M1006 dint_bar EN BR VDD pshort W=2 L=0.15 m=1 mult=1

M1007 VDD dint_bar DOUT VDD pshort W=1.26 L=0.15 m=1 mult=1
M1008 DOUT dint_bar GND GND nshort W=0.65 L=0.15 m=1 mult=1

.ENDS sky130_fd_bd_sram__openram_sense_amp
