* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_fom_serif_nmos
.ends
