VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_cell_fom_serifs
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_cell_fom_serifs ;
  ORIGIN -0.070 0.000 ;
  SIZE 0.905 BY 0.245 ;
END sky130_fd_bd_sram__openram_sp_cell_fom_serifs
END LIBRARY

