# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_wlstrap_p
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_wlstrap_p ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  1.410000 BY  1.580000 ;
  PIN vgnd
    ANTENNADIFFAREA  0.043200 ;
    PORT
      LAYER met1 ;
        POLYGON 1.170000 0.630000 1.195000 0.630000 1.195000 0.605000 ;
        RECT 1.170000 0.630000 1.300000 0.635000 ;
        RECT 1.170000 0.635000 1.355000 0.895000 ;
        RECT 1.170000 0.895000 1.300000 1.315000 ;
        RECT 1.195000 0.605000 1.300000 0.630000 ;
        RECT 1.230000 0.000000 1.300000 0.605000 ;
        RECT 1.230000 1.315000 1.300000 1.580000 ;
    END
    PORT
      LAYER met2 ;
        RECT -0.055000 0.635000 1.355000 0.895000 ;
    END
  END vgnd
  OBS
    LAYER li1 ;
      RECT 0.000000 0.705000 0.085000 0.875000 ;
      RECT 0.280000 0.200000 0.450000 0.370000 ;
      RECT 0.565000 0.160000 0.735000 0.330000 ;
      RECT 0.565000 0.715000 0.735000 0.885000 ;
      RECT 0.565000 1.055000 0.735000 1.225000 ;
      RECT 0.825000 0.605000 0.995000 0.775000 ;
      RECT 0.825000 0.965000 0.995000 1.135000 ;
      RECT 0.850000 0.200000 1.020000 0.370000 ;
      RECT 1.215000 0.705000 1.300000 0.875000 ;
    LAYER met1 ;
      POLYGON  0.105000 0.630000 0.130000 0.630000 0.105000 0.605000 ;
      POLYGON  0.270000 0.570000 0.270000 0.510000 0.210000 0.510000 ;
      POLYGON  0.380000 0.580000 0.510000 0.580000 0.380000 0.450000 ;
      POLYGON  0.520000 0.105000 0.525000 0.105000 0.525000 0.100000 ;
      POLYGON  0.525000 0.100000 0.555000 0.100000 0.555000 0.070000 ;
      POLYGON  0.555000 0.410000 0.555000 0.375000 0.520000 0.375000 ;
      POLYGON  0.745000 0.100000 0.775000 0.100000 0.745000 0.070000 ;
      POLYGON  0.745000 0.410000 0.780000 0.375000 0.745000 0.375000 ;
      POLYGON  0.775000 0.105000 0.780000 0.105000 0.775000 0.100000 ;
      POLYGON  0.790000 0.580000 0.920000 0.580000 0.920000 0.450000 ;
      POLYGON  1.030000 0.570000 1.090000 0.510000 1.030000 0.510000 ;
      RECT -0.055000 0.635000 0.130000 0.895000 ;
      RECT  0.000000 0.000000 0.070000 0.605000 ;
      RECT  0.000000 0.605000 0.105000 0.630000 ;
      RECT  0.000000 0.630000 0.130000 0.635000 ;
      RECT  0.000000 0.895000 0.130000 1.315000 ;
      RECT  0.000000 1.315000 0.070000 1.580000 ;
      RECT  0.210000 0.000000 0.380000 0.510000 ;
      RECT  0.270000 0.510000 0.380000 0.580000 ;
      RECT  0.270000 0.580000 0.510000 1.580000 ;
      RECT  0.520000 0.105000 0.780000 0.375000 ;
      RECT  0.525000 0.100000 0.775000 0.105000 ;
      RECT  0.555000 0.070000 0.745000 0.100000 ;
      RECT  0.555000 0.375000 0.745000 0.410000 ;
      RECT  0.790000 0.580000 1.030000 1.580000 ;
      RECT  0.920000 0.000000 1.090000 0.510000 ;
      RECT  0.920000 0.510000 1.030000 0.580000 ;
    LAYER met2 ;
      RECT 0.000000 0.295000 1.300000 0.465000 ;
      RECT 0.000000 1.065000 1.300000 1.285000 ;
      RECT 0.490000 0.120000 0.810000 0.295000 ;
      RECT 0.520000 0.115000 0.780000 0.120000 ;
    LAYER pwell ;
      RECT 0.415000 0.610000 0.885000 1.260000 ;
    LAYER via ;
      RECT 0.520000 0.115000 0.780000 0.375000 ;
  END
END sky130_fd_bd_sram__sram_sp_wlstrap_p
END LIBRARY
