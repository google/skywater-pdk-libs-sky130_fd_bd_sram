* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell_fom_serifs.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cell_fom_serifs
.ends
