magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1271 1751 1587
<< via1 >>
rect -11 290 26 327
rect 454 132 491 184
rect -11 -11 26 26
<< metal2 >>
rect 26 290 41 316
rect 0 279 41 290
rect 108 244 480 292
rect 108 195 156 244
rect 0 147 156 195
rect 439 184 480 196
rect 439 168 454 184
rect 324 132 454 168
rect 324 120 480 132
rect 324 37 372 120
rect 0 26 372 37
rect 26 0 372 26
<< metal3 >>
rect 0 275 480 316
rect 0 101 480 215
rect 0 0 480 41
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_cell_met23_opt5.gds
string GDS_END 1090
string GDS_START 174
<< end >>
