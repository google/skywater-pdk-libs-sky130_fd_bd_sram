VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_wlstrap_p_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_wlstrap_p_ce ;
  ORIGIN 0.055 0.000 ;
  SIZE 1.410 BY 1.580 ;
  OBS
      LAYER pwell ;
        RECT 0.415 0.610 0.885 1.260 ;
      LAYER li1 ;
        RECT 0.565 1.055 0.735 1.225 ;
        RECT 0.825 0.965 0.995 1.135 ;
        RECT 0.000 0.705 0.085 0.875 ;
        RECT 0.565 0.715 0.735 0.885 ;
        RECT 0.825 0.605 0.995 0.775 ;
        RECT 1.215 0.705 1.300 0.875 ;
        RECT 0.280 0.200 0.450 0.370 ;
        RECT 0.565 0.160 0.735 0.330 ;
        RECT 0.850 0.200 1.020 0.370 ;
      LAYER met1 ;
        RECT 0.000 1.315 0.070 1.580 ;
        RECT 0.000 0.895 0.130 1.315 ;
        RECT -0.055 0.635 0.130 0.895 ;
        RECT 0.000 0.630 0.130 0.635 ;
        RECT 0.000 0.605 0.105 0.630 ;
        POLYGON 0.105 0.630 0.130 0.630 0.105 0.605 ;
        RECT 0.000 0.000 0.070 0.605 ;
        RECT 0.270 0.580 0.510 1.580 ;
        POLYGON 0.270 0.570 0.270 0.510 0.210 0.510 ;
        RECT 0.270 0.510 0.380 0.580 ;
        RECT 0.210 0.000 0.380 0.510 ;
        POLYGON 0.380 0.580 0.510 0.580 0.380 0.450 ;
        RECT 0.790 0.580 1.030 1.580 ;
        RECT 1.230 1.315 1.300 1.580 ;
        RECT 1.170 0.895 1.300 1.315 ;
        RECT 1.170 0.635 1.355 0.895 ;
        RECT 1.170 0.630 1.300 0.635 ;
        POLYGON 1.170 0.630 1.195 0.630 1.195 0.605 ;
        RECT 1.195 0.605 1.300 0.630 ;
        POLYGON 0.790 0.580 0.920 0.580 0.920 0.450 ;
        RECT 0.920 0.510 1.030 0.580 ;
        POLYGON 1.030 0.570 1.090 0.510 1.030 0.510 ;
        POLYGON 0.555 0.410 0.555 0.375 0.520 0.375 ;
        RECT 0.555 0.375 0.745 0.410 ;
        POLYGON 0.745 0.410 0.780 0.375 0.745 0.375 ;
        RECT 0.520 0.105 0.780 0.375 ;
        POLYGON 0.520 0.105 0.525 0.105 0.525 0.100 ;
        RECT 0.525 0.100 0.775 0.105 ;
        POLYGON 0.775 0.105 0.780 0.105 0.775 0.100 ;
        POLYGON 0.525 0.100 0.555 0.100 0.555 0.070 ;
        RECT 0.555 0.070 0.745 0.100 ;
        POLYGON 0.745 0.100 0.775 0.100 0.745 0.070 ;
        RECT 0.920 0.000 1.090 0.510 ;
        RECT 1.230 0.000 1.300 0.605 ;
      LAYER via ;
        RECT 0.520 0.115 0.780 0.375 ;
      LAYER met2 ;
        RECT -0.055 0.635 0.130 0.895 ;
        RECT 1.170 0.635 1.355 0.895 ;
        RECT 0.490 0.120 0.810 0.440 ;
        RECT 0.520 0.115 0.780 0.120 ;
  END
END sky130_fd_bd_sram__sram_sp_wlstrap_p_ce
END LIBRARY

