# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_blkinv_met23
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_blkinv_met23 ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  3.165000 BY  0.900000 ;
  OBS
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000 0.130000 ;
      RECT -0.055000  0.660000 0.130000 0.845000 ;
      RECT  2.925000 -0.055000 3.110000 0.130000 ;
      RECT  2.925000  0.660000 3.110000 0.845000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 -0.040000 ;
      RECT -0.055000 -0.040000 0.140000  0.000000 ;
      RECT -0.055000  0.000000 0.240000  0.130000 ;
      RECT -0.055000  0.660000 0.240000  0.790000 ;
      RECT -0.055000  0.790000 0.140000  0.830000 ;
      RECT -0.055000  0.830000 0.130000  0.845000 ;
      RECT -0.040000  0.130000 0.240000  0.140000 ;
      RECT -0.040000  0.650000 0.240000  0.660000 ;
      RECT  0.000000  0.140000 0.240000  0.650000 ;
      RECT  1.600000  0.000000 3.110000  0.130000 ;
      RECT  1.600000  0.130000 3.055000  0.660000 ;
      RECT  1.600000  0.660000 3.110000  0.790000 ;
      RECT  2.925000 -0.055000 3.110000  0.000000 ;
      RECT  2.925000  0.790000 3.110000  0.845000 ;
    LAYER met3 ;
      RECT -0.040000 -0.040000 0.140000 0.000000 ;
      RECT -0.040000  0.000000 3.055000 0.140000 ;
      RECT -0.040000  0.650000 3.055000 0.790000 ;
      RECT -0.040000  0.790000 0.140000 0.830000 ;
      RECT  0.000000  0.140000 3.055000 0.205000 ;
      RECT  0.000000  0.205000 0.205000 0.585000 ;
      RECT  0.000000  0.585000 3.055000 0.650000 ;
    LAYER via2 ;
      RECT -0.040000 -0.040000 0.140000 0.140000 ;
  END
END sky130_fd_bd_sram__sram_dp_blkinv_met23
END LIBRARY
