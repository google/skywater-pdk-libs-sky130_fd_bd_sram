magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1312 -1237 1227 1552
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optb  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optb_0
timestamp 0
transform 1 0 -52 0 1 23
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optb  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optb_1
timestamp 0
transform 1 0 -52 0 1 261
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta_0
timestamp 0
transform 1 0 -52 0 1 291
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_opta_1
timestamp 0
transform 1 0 -52 0 1 53
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optd  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optd_0
timestamp 0
transform 1 0 -34 0 1 181
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optd  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optd_1
timestamp 0
transform 1 0 -34 0 1 103
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optc  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optc_0
timestamp 0
transform 1 0 -34 0 1 211
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optc  sky130_fd_bd_sram__sram_dp_swldrv_opt1_poly_siz_optc_1
timestamp 0
transform 1 0 -34 0 1 133
box 0 0 1 1
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_swldrv_p1m_siz_a.gds
string GDS_END 1654
string GDS_START 1042
<< end >>
