* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_nand3_dec GND VDD
X0 GND C a_128_208# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VDD C Z VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 Z B VDD VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_128_136# A Z GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VDD A Z VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_128_208# B a_128_136# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
