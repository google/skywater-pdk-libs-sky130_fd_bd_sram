* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell
X0 a_38_54# a_16_24# a_38_0# VSUBS sky130_fd_pr__special_nfet_pass ad=4.375e+10p pd=920000u as=1.68e+10p ps=520000u w=140000u l=150000u
X1 a_38_212# a_16_182# a_0_142# VSUBS sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=8.08e+10p ps=1.28e+06u w=210000u l=150000u
X2 a_38_292# a_16_262# a_38_212# VSUBS sky130_fd_pr__special_nfet_pass ad=1.68e+10p pd=520000u as=4.375e+10p ps=920000u w=140000u l=150000u
X3 a_174_212# a_16_262# a_174_212# w_138_13# sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
X4 a_174_54# a_16_24# a_174_54# w_138_13# sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
X5 a_174_134# a_16_104# a_174_54# w_138_13# sky130_fd_pr__special_pfet_pass ad=6.4e+10p pd=1.14e+06u as=0p ps=0u w=140000u l=150000u
X6 a_174_212# a_16_182# a_174_134# w_138_13# sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X7 a_0_142# a_16_104# a_38_54# VSUBS sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends
