* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_nand2_dec GND VDD
X0 Z A VDD VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VDD B Z VDD sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 a_196_224# B GND GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 Z A a_196_224# GND sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
