# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_dp_nand4_dec
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_dp_nand4_dec ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.610000 BY  1.975000 ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.590000 1.445000 1.920000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.110000 1.085000 1.440000 1.255000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.630000 0.725000 0.960000 0.895000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.365000 0.480000 0.535000 ;
    END
  END D
  PIN GND
    ANTENNADIFFAREA  0.473400 ;
    PORT
      LAYER met1 ;
        RECT 2.270000 -0.305000 2.520000 1.795000 ;
      LAYER pwell ;
        RECT 1.350000 -0.085000 1.760000 0.095000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.324800 ;
    PORT
      LAYER met1 ;
        RECT 4.400000 -0.165000 4.640000 1.765000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.270000 -0.165000 6.510000 1.815000 ;
      LAYER nwell ;
        RECT 3.110000 -0.300000 7.660000 2.660000 ;
    END
  END VDD
  PIN Z
    ANTENNADIFFAREA  0.336000 ;
    PORT
      LAYER li1 ;
        RECT 5.910000 1.405000 7.360000 1.575000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT 1.350000 -0.090000 2.750000 0.100000 ;
      RECT 2.100000  1.585000 3.160000 1.760000 ;
      RECT 2.960000  1.405000 5.200000 1.575000 ;
      RECT 2.960000  1.575000 3.160000 1.585000 ;
      RECT 3.575000  0.470000 4.475000 0.475000 ;
      RECT 3.575000  0.475000 4.690000 0.640000 ;
      RECT 3.575000  0.640000 3.770000 0.950000 ;
      RECT 3.595000  0.950000 3.770000 0.960000 ;
      RECT 3.595000  0.960000 3.765000 1.405000 ;
      RECT 4.350000  0.640000 4.690000 0.645000 ;
      RECT 4.350000  0.935000 4.685000 1.105000 ;
      RECT 5.910000  0.490000 6.345000 0.495000 ;
      RECT 5.910000  0.495000 6.560000 0.660000 ;
      RECT 6.220000  0.660000 6.560000 0.665000 ;
      RECT 6.220000  0.925000 6.555000 1.105000 ;
      RECT 6.300000 -0.165000 6.480000 0.165000 ;
    LAYER mcon ;
      RECT 2.310000 -0.085000 2.480000 0.085000 ;
      RECT 4.435000  0.935000 4.605000 1.105000 ;
      RECT 6.305000  0.930000 6.475000 1.100000 ;
      RECT 6.310000 -0.085000 6.480000 0.085000 ;
  END
END sky130_fd_bd_sram__openram_dp_nand4_dec
END LIBRARY
