# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sense_amp
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sense_amp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.500000 BY  11.28000 ;
  PIN BL
    ANTENNADIFFAREA  0.540000 ;
    PORT
      LAYER met1 ;
        RECT 0.920000 5.420000 1.210000  5.650000 ;
        RECT 0.980000 0.000000 1.150000  5.420000 ;
        RECT 0.980000 5.650000 1.150000 11.280000 ;
    END
  END BL
  PIN BR
    ANTENNADIFFAREA  0.540000 ;
    PORT
      LAYER met1 ;
        RECT 1.360000 0.000000 1.500000  5.420000 ;
        RECT 1.360000 5.420000 1.700000  5.710000 ;
        RECT 1.360000 5.710000 1.500000 11.280000 ;
    END
  END BR
  PIN DOUT
    ANTENNADIFFAREA  0.553900 ;
    PORT
      LAYER met1 ;
        RECT 0.520000 0.000000 0.750000 1.270000 ;
    END
  END DOUT
  PIN E_N
    ANTENNAGATEAREA  0.697500 ;
    PORT
      LAYER met1 ;
        RECT 0.470000 10.820000 0.760000 11.120000 ;
    END
  END E_N
  PIN GND
    ANTENNADIFFAREA  0.266700 ;
    PORT
      LAYER met1 ;
        RECT 1.790000 0.355000 2.020000 0.725000 ;
      LAYER pwell ;
        RECT 1.820000 0.415000 1.990000 0.875000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.140000 10.025000 2.370000 10.395000 ;
      LAYER pwell ;
        RECT 2.170000 10.085000 2.340000 10.545000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.435100 ;
    PORT
      LAYER met1 ;
        RECT 1.690000 6.170000 2.000000 6.510000 ;
      LAYER nwell ;
        RECT -0.800000 1.320000 3.420000 2.620000 ;
        RECT -0.800000 2.620000 3.410000 8.070000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.790000 1.960000 2.020000 2.340000 ;
    END
  END VDD
  OBS
    LAYER li1 ;
      RECT 0.530000 10.880000 1.450000 11.050000 ;
      RECT 0.530000 11.050000 0.700000 11.060000 ;
      RECT 0.540000  3.280000 0.710000  9.150000 ;
      RECT 0.550000  0.300000 0.720000  2.790000 ;
      RECT 0.980000  0.300000 1.160000  0.580000 ;
      RECT 0.980000  0.580000 1.990000  0.760000 ;
      RECT 0.980000  0.760000 1.160000  1.000000 ;
      RECT 0.980000  3.470000 1.150000  5.620000 ;
      RECT 0.980000  6.260000 1.930000  6.430000 ;
      RECT 0.980000  6.430000 1.150000  7.900000 ;
      RECT 0.980000  8.425000 1.150000 10.710000 ;
      RECT 0.990000  1.490000 1.160000  2.060000 ;
      RECT 0.990000  2.060000 1.990000  2.230000 ;
      RECT 0.990000  2.230000 1.160000  2.790000 ;
      RECT 1.420000  6.600000 1.590000  9.415000 ;
      RECT 1.420000  9.415000 1.870000  9.585000 ;
      RECT 1.420000 10.005000 1.590000 10.255000 ;
      RECT 1.420000 10.255000 2.340000 10.425000 ;
      RECT 1.420000 10.425000 1.590000 10.710000 ;
      RECT 1.500000  3.490000 1.670000  5.650000 ;
      RECT 1.760000  6.430000 1.930000  6.570000 ;
      RECT 1.760000  6.570000 2.190000  6.740000 ;
      RECT 1.820000  0.415000 1.990000  0.580000 ;
      RECT 1.820000  0.760000 1.990000  0.835000 ;
      RECT 1.940000  2.740000 2.110000  5.780000 ;
      RECT 1.940000  5.780000 2.370000  5.950000 ;
      RECT 2.100000  5.950000 2.370000  6.110000 ;
      RECT 2.170000 10.085000 2.340000 10.255000 ;
      RECT 2.170000 10.425000 2.340000 10.505000 ;
    LAYER mcon ;
      RECT 0.530000 10.885000 0.700000 11.055000 ;
      RECT 0.550000  1.040000 0.720000  1.210000 ;
      RECT 0.980000  5.450000 1.150000  5.620000 ;
      RECT 1.500000  5.480000 1.670000  5.650000 ;
      RECT 1.760000  6.260000 1.930000  6.430000 ;
      RECT 1.820000  2.060000 1.990000  2.230000 ;
  END
END sky130_fd_bd_sram__openram_sense_amp
END LIBRARY
