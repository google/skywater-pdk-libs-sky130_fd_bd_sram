# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_nand4_dec
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_nand4_dec ;
  ORIGIN  2.375000 -0.175000 ;
  SIZE  9.675000 BY  1.580000 ;
  PIN GND
    ANTENNADIFFAREA  0.389450 ;
    PORT
      LAYER met1 ;
        RECT -1.685000 0.925000 -1.450000 1.465000 ;
      LAYER pwell ;
        RECT -0.295000 1.300000 -0.025000 1.715000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.859175 ;
    PORT
      LAYER met1 ;
        RECT 3.360000 0.070000 3.600000 1.840000 ;
        RECT 5.690000 0.070000 5.930000 1.380000 ;
        RECT 5.690000 1.380000 7.300000 1.620000 ;
        RECT 5.690000 1.620000 5.930000 1.745000 ;
      LAYER nwell ;
        RECT 2.070000 -0.300000 7.325000 2.370000 ;
        RECT 5.430000  2.370000 7.325000 2.375000 ;
    END
  END VDD
  OBS
    LAYER li1 ;
      RECT -2.375000 0.780000 -2.045000 0.950000 ;
      RECT -1.870000 1.005000 -1.210000 1.200000 ;
      RECT -1.865000 0.530000 -1.215000 0.725000 ;
      RECT -1.685000 1.200000 -1.450000 1.580000 ;
      RECT -1.685000 1.580000  0.005000 1.755000 ;
      RECT -0.995000 0.865000 -0.655000 0.950000 ;
      RECT -0.995000 0.950000 -0.570000 1.160000 ;
      RECT -0.350000 0.880000 -0.020000 1.050000 ;
      RECT -0.295000 1.340000  0.005000 1.580000 ;
      RECT  0.200000 0.430000  0.530000 0.600000 ;
      RECT  0.200000 1.330000  0.530000 1.500000 ;
      RECT  0.700000 1.455000  1.360000 1.650000 ;
      RECT  0.710000 0.305000  6.780000 0.475000 ;
      RECT  1.630000 1.215000  1.970000 1.300000 ;
      RECT  1.630000 1.300000  2.055000 1.510000 ;
      RECT  2.555000 0.475000  2.725000 1.275000 ;
      RECT  2.555000 1.275000  3.650000 1.440000 ;
      RECT  2.555000 1.440000  3.435000 1.445000 ;
      RECT  3.310000 0.770000  5.975000 0.940000 ;
      RECT  3.310000 1.270000  3.650000 1.275000 ;
      RECT  4.610000 1.215000  4.950000 1.300000 ;
      RECT  4.610000 1.300000  5.035000 1.510000 ;
      RECT  5.645000 1.255000  6.315000 1.425000 ;
      RECT  6.145000 0.475000  6.315000 1.255000 ;
      RECT  6.675000 0.715000  7.015000 1.010000 ;
      RECT  6.820000 1.400000  7.150000 1.590000 ;
    LAYER mcon ;
      RECT -1.650000 0.540000 -1.480000 0.710000 ;
      RECT -1.650000 1.015000 -1.480000 1.185000 ;
      RECT -0.915000 0.925000 -0.745000 1.095000 ;
      RECT  0.955000 1.465000  1.125000 1.635000 ;
      RECT  1.710000 1.275000  1.880000 1.445000 ;
      RECT  3.395000 0.770000  3.565000 0.940000 ;
      RECT  4.690000 1.275000  4.860000 1.445000 ;
      RECT  5.725000 0.770000  5.895000 0.940000 ;
      RECT  6.755000 0.775000  6.925000 0.945000 ;
      RECT  6.900000 1.415000  7.070000 1.585000 ;
    LAYER met1 ;
      RECT -1.715000 0.500000  1.385000 0.640000 ;
      RECT -1.715000 0.640000 -1.250000 0.755000 ;
      RECT -0.995000 0.785000 -0.650000 1.100000 ;
      RECT -0.995000 1.100000 -0.655000 1.160000 ;
      RECT  0.895000 0.640000  1.185000 1.700000 ;
      RECT  1.630000 1.135000  1.975000 1.450000 ;
      RECT  1.630000 1.450000  1.970000 1.510000 ;
      RECT  4.610000 1.135000  4.955000 1.450000 ;
      RECT  4.610000 1.450000  4.950000 1.510000 ;
      RECT  6.675000 0.635000  7.015000 1.010000 ;
    LAYER met2 ;
      RECT -0.995000 0.785000 -0.650000 0.855000 ;
      RECT -0.995000 0.855000  7.015000 0.995000 ;
      RECT -0.995000 0.995000 -0.650000 1.090000 ;
      RECT  1.630000 1.135000  1.975000 1.300000 ;
      RECT  1.630000 1.300000  5.045000 1.440000 ;
      RECT  4.610000 1.135000  4.955000 1.300000 ;
      RECT  6.675000 0.635000  7.015000 0.855000 ;
    LAYER via ;
      RECT -0.955000 0.820000 -0.695000 1.080000 ;
      RECT  1.670000 1.170000  1.930000 1.430000 ;
      RECT  4.650000 1.170000  4.910000 1.430000 ;
      RECT  6.715000 0.670000  6.975000 0.930000 ;
  END
END sky130_fd_bd_sram__openram_nand4_dec
END LIBRARY
