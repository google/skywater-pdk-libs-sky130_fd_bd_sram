* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_dp_cell_replica BL0 BL1 BR0 BR1 GND VDD WL0 WL1
X0 a_38_133# VDD GND GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X1 BL1 GND BL1 GND sky130_fd_pr__special_nfet_pass w=105000u l=185000u
X2 a_38_133# WL1 BL1 GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X3 BR0 WL0 VDD GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X4 a_38_n79# GND a_38_n79# GND sky130_fd_pr__special_nfet_pass w=105000u l=185000u
X5 a_400_n79# GND a_400_n79# GND sky130_fd_pr__special_nfet_pass w=105000u l=185000u
X6 BR1 GND BR1 GND sky130_fd_pr__special_nfet_pass w=105000u l=185000u
X7 GND a_38_133# VDD GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X8 VDD a_38_133# GND GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X9 BL0 WL0 a_38_133# GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X10 VDD WL1 BR1 GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
X11 GND VDD a_38_133# GND sky130_fd_pr__special_nfet_latch w=210000u l=150000u
.ends
