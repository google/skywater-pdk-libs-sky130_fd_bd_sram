
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.SUBCKT sky130_fd_bd_sram__openram_cell_1rw_1r_dummy bl0 br0 bl1 br1 wl0 wl1 vdd gnd
** N=14 EP=6 IP=0 FDC=16
*.SEEDPROM

* Bitcell Core
X1 1 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X2 1 wl1 bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X3 2 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X4 2 wl1 br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X5 3 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X6 3 wl0 bl0 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X7 4 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15
X8 4 wl0 br0 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15

* drainOnly NMOS
X9 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08
X10 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08

.ENDS
