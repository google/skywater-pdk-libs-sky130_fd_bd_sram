VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colend
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colend ;
  ORIGIN 0.055 0.000 ;
  SIZE 1.310 BY 2.055 ;
  PIN BL0
    PORT
      LAYER met1 ;
        RECT 0.710 1.595 0.890 2.055 ;
        RECT 0.710 0.000 0.850 1.595 ;
        POLYGON 0.850 1.595 0.890 1.595 0.850 1.555 ;
    END
  END BL0
  PIN BL1
    ANTENNADIFFAREA 0.016800 ;
    PORT
      LAYER li1 ;
        RECT 0.335 0.075 0.505 0.085 ;
        RECT 0.870 0.075 1.010 0.085 ;
        RECT 0.070 0.000 1.130 0.075 ;
      LAYER mcon ;
        RECT 0.335 0.000 0.505 0.085 ;
      LAYER met1 ;
        RECT 0.305 1.590 0.485 2.055 ;
        POLYGON 0.305 1.590 0.345 1.590 0.345 1.550 ;
        RECT 0.345 0.145 0.485 1.590 ;
        RECT 0.300 0.000 0.540 0.145 ;
    END
  END BL1
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.050 1.955 1.200 2.055 ;
        RECT 1.050 1.695 1.255 1.955 ;
        RECT 1.050 1.595 1.200 1.695 ;
        POLYGON 1.050 1.595 1.130 1.595 1.130 1.515 ;
        RECT 1.130 0.000 1.200 1.595 ;
      LAYER via ;
        RECT 1.070 1.695 1.255 1.955 ;
      LAYER met2 ;
        RECT 0.000 1.955 1.200 2.055 ;
        RECT 0.000 1.695 1.255 1.955 ;
        RECT 0.000 1.600 1.200 1.695 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 1.025 0.090 2.055 ;
        POLYGON 0.090 1.105 0.170 1.025 0.090 1.025 ;
        RECT 0.000 1.005 0.170 1.025 ;
        RECT -0.055 0.745 0.170 1.005 ;
        RECT 0.000 0.730 0.170 0.745 ;
        RECT 0.000 0.000 0.070 0.730 ;
        POLYGON 0.070 0.730 0.170 0.730 0.070 0.630 ;
      LAYER met2 ;
        RECT 0.000 1.005 1.200 1.030 ;
        RECT -0.055 0.745 1.200 1.005 ;
        RECT 0.000 0.580 1.200 0.745 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 0.000 0.480 2.055 ;
      LAYER pwell ;
        RECT 0.700 0.530 1.200 1.680 ;
      LAYER li1 ;
        RECT 0.000 1.175 1.200 1.875 ;
        RECT 0.000 0.990 0.340 1.175 ;
        RECT 0.520 0.810 1.200 1.005 ;
        RECT 0.000 0.275 1.200 0.810 ;
      LAYER met2 ;
        RECT 0.000 1.180 1.200 1.460 ;
        RECT 0.000 0.020 1.200 0.405 ;
  END
END sky130_fd_bd_sram__sram_sp_colend
END LIBRARY

