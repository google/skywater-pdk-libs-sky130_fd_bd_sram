* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_write_driver" ******************************

.SUBCKT sky130_fd_bd_sram__openram_write_driver DIN BL BR EN VDD GND

**** Inverter to conver Data_in to data_in_bar ******
* din_bar = inv(DIN)
M_1 din_bar DIN GND GND nshort W=0.36 L=0.15 m=1 mult=1
M_2 din_bar DIN VDD VDD pshort W=0.55 L=0.15 m=1 mult=1

**** 2input nand gate follwed by inverter to drive BL ******
* din_bar_gated = nand(EN, DIN)
M_3 din_bar_gated EN net_7 GND nshort W=0.55 L=0.15 m=1 mult=1
M_4 net_7 DIN GND GND nshort W=0.55 L=0.15 m=1 mult=1
M_5 din_bar_gated EN VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
M_6 din_bar_gated DIN VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
* din_bar_gated_bar = inv(din_bar_gated)
M_7 din_bar_gated_bar din_bar_gated VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
M_8 din_bar_gated_bar din_bar_gated GND GND nshort W=0.36 L=0.15 m=1 mult=1

**** 2input nand gate follwed by inverter to drive BR******
* din_gated = nand(EN, din_bar)
M_9 din_gated EN VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
M_10 din_gated EN net_8 GND nshort W=0.55 L=0.15 m=1 mult=1
M_11 net_8 din_bar GND GND nshort W=0.55 L=0.15 m=1 mult=1
M_12 din_gated din_bar VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
* din_gated_bar = inv(din_gated)
M_13 din_gated_bar din_gated VDD VDD pshort W=0.55 L=0.15 m=1 mult=1
M_14 din_gated_bar din_gated GND GND nshort W=0.36 L=0.15 m=1 mult=1

************************************************
* pull down with EN enable
M_15 BL din_gated_bar GND GND nshort W=1 L=0.15 m=1 mult=1
M_16 BR din_bar_gated_bar GND GND nshort W=1 L=0.15 m=1 mult=1

.ENDS sky130_fd_bd_sram__openram_write_driver
