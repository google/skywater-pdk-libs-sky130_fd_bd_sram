# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sram_dff
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sram_dff ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.840000 BY  7.070000 ;
  PIN CLK
    ANTENNAGATEAREA  1.800000 ;
    PORT
      LAYER met2 ;
        RECT 1.845000 3.460000 2.115000 3.780000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.600000 ;
    PORT
      LAYER met2 ;
        RECT 0.685000 2.690000 1.015000 2.950000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.060000 ;
    ANTENNAGATEAREA  0.600000 ;
    PORT
      LAYER met2 ;
        RECT 5.410000 3.045000 5.740000 3.305000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  1.800000 ;
    ANTENNAGATEAREA  0.600000 ;
    PORT
      LAYER met2 ;
        RECT 5.020000 2.290000 5.350000 2.550000 ;
    END
  END Q_N
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.100000 5.840000 0.100000 ;
      RECT 0.000000  6.980000 5.840000 7.160000 ;
      RECT 0.180000  0.510000 0.350000 1.350000 ;
      RECT 0.180000  2.335000 1.365000 2.505000 ;
      RECT 0.180000  3.935000 0.350000 6.560000 ;
      RECT 0.205000  3.135000 0.735000 3.305000 ;
      RECT 0.205000  3.535000 5.660000 3.705000 ;
      RECT 0.610000  0.100000 0.780000 1.350000 ;
      RECT 0.610000  4.020000 0.780000 6.980000 ;
      RECT 0.685000  2.735000 1.015000 2.905000 ;
      RECT 1.195000  2.505000 1.365000 2.660000 ;
      RECT 1.195000  2.660000 2.530000 2.830000 ;
      RECT 1.245000  3.030000 1.415000 3.535000 ;
      RECT 1.400000  0.510000 1.740000 1.350000 ;
      RECT 1.400000  4.020000 1.740000 6.560000 ;
      RECT 1.485000  3.935000 1.655000 4.020000 ;
      RECT 1.640000  1.935000 2.065000 2.105000 ;
      RECT 2.280000  1.935000 2.610000 2.105000 ;
      RECT 2.280000  3.115000 2.610000 3.285000 ;
      RECT 2.360000  0.100000 2.530000 1.350000 ;
      RECT 2.360000  2.105000 2.530000 2.660000 ;
      RECT 2.360000  2.830000 2.530000 3.115000 ;
      RECT 2.360000  4.020000 2.530000 6.980000 ;
      RECT 2.915000  1.935000 3.245000 2.105000 ;
      RECT 2.995000  2.105000 3.165000 3.535000 ;
      RECT 3.150000  0.510000 3.490000 1.350000 ;
      RECT 3.150000  4.020000 3.490000 6.560000 ;
      RECT 3.235000  1.350000 3.405000 1.535000 ;
      RECT 3.235000  1.535000 5.230000 1.705000 ;
      RECT 3.235000  3.935000 3.405000 4.020000 ;
      RECT 3.395000  2.335000 4.710000 2.505000 ;
      RECT 3.475000  3.030000 3.645000 3.535000 ;
      RECT 3.875000  2.735000 5.660000 2.905000 ;
      RECT 4.110000  0.100000 4.280000 1.350000 ;
      RECT 4.110000  4.020000 4.280000 6.980000 ;
      RECT 4.390000  3.135000 4.720000 3.305000 ;
      RECT 4.470000  3.305000 4.640000 3.535000 ;
      RECT 4.540000  0.510000 4.710000 1.355000 ;
      RECT 4.540000  3.935000 4.710000 6.560000 ;
      RECT 5.060000  0.100000 5.230000 1.350000 ;
      RECT 5.060000  1.705000 5.230000 2.335000 ;
      RECT 5.060000  2.335000 5.465000 2.505000 ;
      RECT 5.060000  4.020000 5.230000 6.980000 ;
      RECT 5.490000  0.510000 5.660000 1.355000 ;
      RECT 5.490000  2.905000 5.660000 3.260000 ;
      RECT 5.490000  3.935000 5.660000 6.560000 ;
    LAYER mcon ;
      RECT 0.180000 1.135000 0.350000 1.305000 ;
      RECT 0.565000 3.135000 0.735000 3.305000 ;
      RECT 0.765000 2.735000 0.935000 2.905000 ;
      RECT 1.485000 1.135000 1.655000 1.305000 ;
      RECT 1.895000 1.935000 2.065000 2.105000 ;
      RECT 1.895000 3.535000 2.065000 3.705000 ;
      RECT 3.235000 1.135000 3.405000 1.305000 ;
      RECT 4.540000 1.135000 4.710000 1.305000 ;
      RECT 4.540000 2.335000 4.710000 2.505000 ;
      RECT 5.100000 2.335000 5.270000 2.505000 ;
      RECT 5.490000 1.135000 5.660000 1.305000 ;
      RECT 5.490000 3.090000 5.660000 3.260000 ;
    LAYER met1 ;
      RECT 0.120000 1.105000 0.410000 1.335000 ;
      RECT 0.120000 2.305000 0.410000 2.535000 ;
      RECT 0.120000 3.905000 0.410000 4.135000 ;
      RECT 0.180000 1.335000 0.350000 2.305000 ;
      RECT 0.180000 2.535000 0.350000 3.905000 ;
      RECT 0.505000 3.105000 0.795000 3.135000 ;
      RECT 0.505000 3.135000 1.655000 3.305000 ;
      RECT 0.505000 3.305000 0.795000 3.335000 ;
      RECT 0.685000 2.690000 1.015000 2.950000 ;
      RECT 1.425000 1.105000 1.715000 1.335000 ;
      RECT 1.425000 3.905000 1.715000 4.135000 ;
      RECT 1.485000 1.335000 1.655000 3.135000 ;
      RECT 1.485000 3.305000 1.655000 3.905000 ;
      RECT 1.835000 1.905000 2.125000 2.135000 ;
      RECT 1.835000 3.505000 2.125000 3.735000 ;
      RECT 1.845000 1.860000 2.115000 1.905000 ;
      RECT 1.845000 2.135000 2.115000 2.180000 ;
      RECT 1.845000 3.460000 2.115000 3.505000 ;
      RECT 1.845000 3.735000 2.115000 3.780000 ;
      RECT 1.895000 2.180000 2.065000 3.460000 ;
      RECT 3.175000 1.105000 3.465000 1.335000 ;
      RECT 3.175000 3.905000 3.465000 4.135000 ;
      RECT 3.235000 1.335000 3.405000 3.905000 ;
      RECT 4.480000 1.105000 4.770000 1.335000 ;
      RECT 4.480000 2.305000 4.770000 2.535000 ;
      RECT 4.480000 3.905000 4.770000 4.135000 ;
      RECT 4.540000 1.335000 4.710000 2.305000 ;
      RECT 4.540000 2.535000 4.710000 3.905000 ;
      RECT 5.020000 2.290000 5.350000 2.550000 ;
      RECT 5.410000 3.045000 5.740000 3.305000 ;
      RECT 5.430000 1.105000 5.720000 1.335000 ;
      RECT 5.430000 3.905000 5.720000 4.135000 ;
      RECT 5.490000 1.335000 5.660000 3.045000 ;
      RECT 5.490000 3.305000 5.660000 3.905000 ;
    LAYER nwell ;
      RECT -0.040000 3.380000 5.880000 7.335000 ;
    LAYER pwell ;
      RECT 0.140000 -0.085000 0.550000 0.085000 ;
      RECT 0.820000 -0.085000 1.230000 0.085000 ;
      RECT 1.500000 -0.085000 1.910000 0.085000 ;
      RECT 2.180000 -0.085000 2.590000 0.085000 ;
      RECT 2.860000 -0.085000 3.270000 0.085000 ;
      RECT 3.540000 -0.085000 3.950000 0.085000 ;
      RECT 4.220000 -0.085000 4.630000 0.085000 ;
      RECT 4.900000 -0.085000 5.310000 0.085000 ;
    LAYER via ;
      RECT 0.720000 2.690000 0.980000 2.950000 ;
      RECT 1.850000 3.490000 2.110000 3.750000 ;
      RECT 5.055000 2.290000 5.315000 2.550000 ;
      RECT 5.445000 3.045000 5.705000 3.305000 ;
  END
END sky130_fd_bd_sram__openram_sram_dff
END LIBRARY
