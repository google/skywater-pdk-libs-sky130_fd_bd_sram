magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1261 1261 1261
use sky130_fd_bd_sram__sram_dp_licon_05  sky130_fd_bd_sram__sram_dp_licon_05_0
timestamp 0
transform 1 0 0 0 -1 0
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_licon_05  sky130_fd_bd_sram__sram_dp_licon_05_1
timestamp 0
transform 1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_licon_1.gds
string GDS_END 424
string GDS_START 294
<< end >>
