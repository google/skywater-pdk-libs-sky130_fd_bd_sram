# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_base
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_base ;
  ORIGIN  3.055000  0.000000 ;
  SIZE  3.055000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT -3.055000 0.000000 -2.740000 0.410000 ;
      RECT -2.545000 0.090000 -1.620000 0.405000 ;
      RECT -2.515000 0.630000 -1.560000 0.685000 ;
      RECT -2.515000 0.685000 -0.265000 0.895000 ;
      RECT -1.575000 1.075000 -0.900000 1.395000 ;
      RECT -0.760000 0.000000 -0.420000 0.160000 ;
      RECT -0.760000 0.160000 -0.565000 0.535000 ;
      RECT -0.760000 1.045000 -0.565000 1.420000 ;
      RECT -0.760000 1.420000 -0.420000 1.580000 ;
      RECT -0.425000 0.320000 -0.070000 0.465000 ;
      RECT -0.425000 0.465000 -0.265000 0.685000 ;
      RECT -0.425000 0.895000 -0.265000 1.115000 ;
      RECT -0.425000 1.115000 -0.070000 1.260000 ;
      RECT -0.275000 0.090000 -0.070000 0.320000 ;
      RECT -0.275000 1.260000 -0.070000 1.490000 ;
      RECT -0.125000 0.625000  0.000000 0.955000 ;
    LAYER mcon ;
      RECT -0.590000 0.000000 -0.420000 0.085000 ;
      RECT -0.590000 1.495000 -0.420000 1.580000 ;
      RECT -0.565000 0.705000 -0.395000 0.875000 ;
      RECT -0.085000 0.705000  0.000000 0.875000 ;
    LAYER met1 ;
      RECT -2.465000 0.000000 -2.215000 1.580000 ;
      RECT -2.015000 0.000000 -1.765000 1.580000 ;
      RECT -1.565000 0.000000 -1.315000 1.580000 ;
      RECT -1.115000 0.000000 -0.865000 1.580000 ;
      RECT -0.685000 0.560000 -0.265000 0.980000 ;
      RECT -0.680000 0.980000 -0.265000 1.045000 ;
      RECT -0.620000 0.000000  0.000000 0.380000 ;
      RECT -0.620000 1.225000  0.000000 1.580000 ;
      RECT -0.085000 0.380000  0.000000 1.225000 ;
    LAYER nwell ;
      RECT -3.055000 0.000000 -1.300000 1.580000 ;
    LAYER pwell ;
      RECT -0.960000 0.000000 -0.460000 0.200000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_base
END LIBRARY
