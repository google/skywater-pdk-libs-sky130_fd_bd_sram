# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_colend_cent_base
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_colend_cent_base ;
  ORIGIN  0.360000  0.000000 ;
  SIZE  1.230000 BY  1.925000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.585000 0.510000 1.925000 ;
      RECT 0.070000 0.090000 0.440000 0.405000 ;
    LAYER mcon ;
      RECT 0.000000 0.775000 0.085000 0.945000 ;
      RECT 0.070000 0.195000 0.240000 0.365000 ;
      RECT 0.425000 0.775000 0.510000 0.945000 ;
    LAYER met1 ;
      RECT -0.135000 0.145000 0.510000 0.405000 ;
      RECT -0.055000 0.730000 0.565000 0.990000 ;
      RECT  0.000000 0.090000 0.510000 0.145000 ;
      RECT  0.000000 0.405000 0.510000 0.730000 ;
      RECT  0.000000 0.990000 0.510000 1.925000 ;
      RECT  0.435000 0.000000 0.510000 0.090000 ;
    LAYER met2 ;
      RECT -0.360000 1.470000 0.870000 1.925000 ;
      RECT -0.135000 0.145000 0.510000 0.405000 ;
      RECT -0.055000 0.730000 0.565000 0.990000 ;
      RECT  0.000000 0.120000 0.510000 0.145000 ;
      RECT  0.000000 0.405000 0.510000 0.730000 ;
      RECT  0.000000 0.990000 0.510000 1.085000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 0.510000 0.205000 ;
    LAYER pwell ;
      RECT 0.000000 0.715000 0.510000 1.795000 ;
    LAYER via ;
      RECT 0.380000 0.730000 0.565000 0.990000 ;
  END
END sky130_fd_bd_sram__sram_dp_colend_cent_base
END LIBRARY
