VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell_addpoly_sizing
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell_addpoly_sizing ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END sky130_fd_bd_sram__sram_sp_cell_addpoly_sizing
END LIBRARY

