magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1277 -1277 1277 1277
use sky130_fd_bd_sram__sram_dp_mcon_05  sky130_fd_bd_sram__sram_dp_mcon_05_0
timestamp 0
transform 1 0 0 0 -1 0
box -17 0 17 17
use sky130_fd_bd_sram__sram_dp_mcon_05  sky130_fd_bd_sram__sram_dp_mcon_05_1
timestamp 0
transform 1 0 0 0 1 0
box -17 0 17 17
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_mcon_1.gds
string GDS_END 418
string GDS_START 292
<< end >>
