VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_rowend_p1m_siz
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_rowend_p1m_siz ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END sky130_fd_bd_sram__sram_sp_rowend_p1m_siz
END LIBRARY

