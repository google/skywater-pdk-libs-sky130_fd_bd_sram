* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrap_p_met2.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrap_p_met2
.ends
