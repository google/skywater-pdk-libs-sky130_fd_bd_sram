# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_cell_half_limcon_optb
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_cell_half_limcon_optb ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.200000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.625000 0.070000 0.955000 ;
      RECT 0.070000 0.000000 0.590000 0.125000 ;
      RECT 0.070000 0.295000 1.200000 0.470000 ;
      RECT 0.070000 1.505000 1.200000 1.580000 ;
      RECT 0.210000 0.470000 1.200000 0.475000 ;
      RECT 0.210000 0.475000 0.380000 1.365000 ;
      RECT 0.490000 1.455000 1.200000 1.505000 ;
      RECT 0.535000 0.670000 0.705000 1.105000 ;
      RECT 0.535000 1.105000 1.200000 1.285000 ;
      RECT 0.730000 0.000000 1.200000 0.125000 ;
      RECT 0.860000 0.655000 1.200000 0.925000 ;
    LAYER mcon ;
      RECT 0.395000 0.000000 0.565000 0.085000 ;
      RECT 0.755000 0.000000 0.925000 0.085000 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
    LAYER met1 ;
      RECT 0.395000 0.000000 0.565000 0.085000 ;
      RECT 0.755000 0.000000 0.925000 0.085000 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
  END
END sky130_fd_bd_sram__sram_dp_cell_half_limcon_optb
END LIBRARY
