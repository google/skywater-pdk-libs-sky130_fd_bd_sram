# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colenda_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colenda_ce ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.200000 BY  2.055000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.275000 1.200000 0.810000 ;
      RECT 0.000000 0.990000 0.340000 1.175000 ;
      RECT 0.000000 1.175000 1.200000 1.875000 ;
      RECT 0.070000 0.000000 1.130000 0.075000 ;
      RECT 0.335000 0.075000 0.505000 0.085000 ;
      RECT 0.520000 0.810000 1.200000 1.005000 ;
    LAYER mcon ;
      RECT 0.335000 0.000000 0.505000 0.085000 ;
    LAYER met1 ;
      POLYGON 0.070000 0.730000 0.170000 0.730000 0.070000 0.630000 ;
      POLYGON 0.090000 1.105000 0.170000 1.025000 0.090000 1.025000 ;
      POLYGON 0.305000 1.590000 0.345000 1.590000 0.345000 1.550000 ;
      POLYGON 0.850000 1.595000 0.890000 1.595000 0.850000 1.555000 ;
      POLYGON 1.050000 1.595000 1.090000 1.595000 1.090000 1.555000 ;
      POLYGON 1.090000 1.555000 1.130000 1.555000 1.130000 1.515000 ;
      RECT 0.000000 0.000000 0.070000 0.730000 ;
      RECT 0.000000 0.730000 0.170000 1.025000 ;
      RECT 0.000000 1.025000 0.090000 2.055000 ;
      RECT 0.300000 0.000000 0.540000 0.145000 ;
      RECT 0.305000 1.590000 0.485000 2.055000 ;
      RECT 0.345000 0.145000 0.485000 1.590000 ;
      RECT 0.710000 0.000000 0.850000 1.595000 ;
      RECT 0.710000 1.595000 0.890000 2.055000 ;
      RECT 1.050000 1.595000 1.200000 2.055000 ;
      RECT 1.090000 1.555000 1.200000 1.595000 ;
      RECT 1.130000 0.000000 1.200000 1.555000 ;
    LAYER nwell ;
      RECT 0.000000 0.000000 0.480000 2.055000 ;
    LAYER pwell ;
      RECT 0.700000 0.530000 1.200000 1.680000 ;
  END
END sky130_fd_bd_sram__sram_sp_colenda_ce
END LIBRARY
