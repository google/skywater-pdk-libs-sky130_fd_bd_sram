# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_swldrv_tap_b
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_swldrv_tap_b ;
  ORIGIN  0.000000  0.895000 ;
  SIZE  2.405000 BY  0.895000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.895000 0.290000 -0.545000 ;
      RECT 0.090000 -0.365000 1.300000 -0.195000 ;
      RECT 0.090000 -0.195000 0.260000 -0.125000 ;
      RECT 0.580000 -0.465000 1.300000 -0.365000 ;
    LAYER mcon ;
      RECT 0.000000 -0.795000 0.085000 -0.625000 ;
    LAYER met1 ;
      RECT 0.000000 -0.795000 0.085000 -0.625000 ;
    LAYER pwell ;
      RECT 0.000000 -0.895000 0.200000 -0.425000 ;
      RECT 0.000000 -0.425000 1.430000 -0.235000 ;
      RECT 0.500000 -0.235000 1.430000 -0.090000 ;
  END
END sky130_fd_bd_sram__sram_dp_swldrv_tap_b
END LIBRARY
