# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_wlstrap
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_wlstrap ;
  ORIGIN  0.150000  0.000000 ;
  SIZE  0.815000 BY  1.580000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.710000 0.085000 0.870000 ;
      RECT 0.070000 0.090000 0.440000 0.405000 ;
      RECT 0.070000 1.175000 0.440000 1.490000 ;
      RECT 0.425000 0.710000 0.615000 0.870000 ;
      RECT 0.445000 0.705000 0.615000 0.710000 ;
      RECT 0.445000 0.870000 0.615000 0.875000 ;
    LAYER mcon ;
      RECT 0.070000 0.195000 0.240000 0.365000 ;
      RECT 0.070000 1.215000 0.240000 1.385000 ;
    LAYER met1 ;
      POLYGON  0.175000 0.500000 0.255000 0.420000 0.175000 0.420000 ;
      POLYGON  0.175000 1.160000 0.255000 1.160000 0.175000 1.080000 ;
      RECT -0.135000 0.145000 0.255000 0.405000 ;
      RECT -0.135000 1.175000 0.255000 1.435000 ;
      RECT  0.000000 0.090000 0.255000 0.145000 ;
      RECT  0.000000 0.405000 0.255000 0.420000 ;
      RECT  0.000000 0.420000 0.175000 0.500000 ;
      RECT  0.000000 1.080000 0.175000 1.160000 ;
      RECT  0.000000 1.160000 0.255000 1.175000 ;
      RECT  0.000000 1.435000 0.255000 1.490000 ;
      RECT  0.350000 0.585000 0.510000 0.660000 ;
      RECT  0.350000 0.660000 0.665000 0.920000 ;
      RECT  0.350000 0.920000 0.510000 0.995000 ;
      RECT  0.435000 0.000000 0.510000 0.585000 ;
      RECT  0.435000 0.995000 0.510000 1.580000 ;
    LAYER met2 ;
      RECT -0.135000 0.145000 0.510000 0.360000 ;
      RECT -0.135000 0.360000 0.200000 0.405000 ;
      RECT -0.135000 1.175000 0.200000 1.220000 ;
      RECT -0.135000 1.220000 0.510000 1.435000 ;
      RECT  0.000000 0.120000 0.510000 0.145000 ;
      RECT  0.000000 0.405000 0.200000 0.430000 ;
      RECT  0.000000 0.670000 0.665000 0.910000 ;
      RECT  0.000000 1.150000 0.200000 1.175000 ;
      RECT  0.000000 1.435000 0.510000 1.460000 ;
      RECT  0.370000 0.600000 0.510000 0.660000 ;
      RECT  0.370000 0.660000 0.665000 0.670000 ;
      RECT  0.370000 0.910000 0.665000 0.920000 ;
      RECT  0.370000 0.920000 0.510000 0.980000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 0.510000 0.205000 ;
      RECT 0.000000 0.505000 0.510000 1.075000 ;
      RECT 0.000000 1.375000 0.510000 1.580000 ;
    LAYER via ;
      RECT 0.405000 0.660000 0.665000 0.920000 ;
  END
END sky130_fd_bd_sram__sram_dp_wlstrap
END LIBRARY
