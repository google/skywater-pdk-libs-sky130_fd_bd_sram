VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_wlstrap_met2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_wlstrap_met2 ;
  ORIGIN 0.000 -0.120 ;
  SIZE 1.300 BY 1.165 ;
  OBS
      LAYER met2 ;
        RECT 0.000 1.025 1.300 1.285 ;
        RECT 0.000 0.635 1.300 0.855 ;
        RECT 0.000 0.295 1.300 0.465 ;
        RECT 0.520 0.120 0.780 0.295 ;
  END
END sky130_fd_bd_sram__sram_sp_wlstrap_met2
END LIBRARY

