# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_colend_half_met23_optb
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_colend_half_met23_optb ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  1.255000 BY  1.980000 ;
  OBS
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000 0.130000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 1.200000 0.130000 ;
      RECT  0.000000  0.130000 1.200000 1.085000 ;
      RECT  0.000000  1.470000 1.200000 1.925000 ;
  END
END sky130_fd_bd_sram__sram_dp_colend_half_met23_optb
END LIBRARY
