VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colenda_cent
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colenda_cent ;
  ORIGIN 0.055 0.000 ;
  SIZE 1.410 BY 2.055 ;
  PIN VNB
    PORT
      LAYER li1 ;
        RECT 0.000 0.275 1.300 0.810 ;
        RECT 0.135 0.015 1.200 0.275 ;
      LAYER mcon ;
        RECT 0.790 0.640 0.960 0.810 ;
        RECT 0.790 0.280 0.960 0.450 ;
      LAYER met1 ;
        RECT 0.750 1.155 1.050 2.055 ;
        RECT 0.750 0.395 0.990 1.155 ;
        POLYGON 0.990 1.155 1.050 1.155 0.990 1.095 ;
        POLYGON 0.990 0.480 1.075 0.395 0.990 0.395 ;
        RECT 0.750 0.380 1.075 0.395 ;
        POLYGON 1.075 0.395 1.090 0.380 1.075 0.380 ;
        RECT 0.750 0.170 1.090 0.380 ;
        POLYGON 0.750 0.170 0.785 0.170 0.785 0.135 ;
        RECT 0.785 0.135 1.090 0.170 ;
        POLYGON 0.785 0.135 0.920 0.135 0.920 0.000 ;
        RECT 0.920 0.000 1.090 0.135 ;
      LAYER via ;
        RECT 0.800 0.135 1.060 0.395 ;
      LAYER met2 ;
        RECT 0.000 0.020 1.300 0.405 ;
    END
  END VNB
  PIN VPB
    ANTENNADIFFAREA 2.034500 ;
    PORT
      LAYER nwell ;
        RECT 0.000 0.000 1.300 2.055 ;
      LAYER li1 ;
        RECT 0.000 0.990 1.300 1.875 ;
      LAYER mcon ;
        RECT 0.295 1.705 0.465 1.875 ;
        RECT 0.295 1.345 0.465 1.515 ;
      LAYER met1 ;
        RECT 0.250 1.155 0.550 2.055 ;
        POLYGON 0.250 1.155 0.310 1.155 0.310 1.095 ;
        POLYGON 0.310 0.480 0.310 0.380 0.210 0.380 ;
        RECT 0.310 0.380 0.550 1.155 ;
        RECT 0.210 0.170 0.550 0.380 ;
        RECT 0.210 0.000 0.380 0.170 ;
        POLYGON 0.380 0.170 0.550 0.170 0.380 0.000 ;
      LAYER via ;
        RECT 0.270 1.190 0.530 1.450 ;
      LAYER met2 ;
        RECT 0.000 1.180 1.300 1.460 ;
    END
  END VPB
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 1.020 0.090 2.055 ;
        POLYGON 1.210 1.105 1.210 1.100 1.205 1.100 ;
        RECT 1.210 1.100 1.300 2.055 ;
        POLYGON 0.090 1.100 0.170 1.020 0.090 1.020 ;
        RECT 0.000 1.005 0.170 1.020 ;
        RECT -0.055 0.745 0.170 1.005 ;
        RECT 0.000 0.730 0.170 0.745 ;
        RECT 0.000 0.000 0.070 0.730 ;
        POLYGON 0.070 0.730 0.170 0.730 0.070 0.630 ;
        POLYGON 1.205 1.100 1.205 1.025 1.130 1.025 ;
        RECT 1.205 1.025 1.300 1.100 ;
        RECT 1.130 1.005 1.300 1.025 ;
        RECT 1.130 0.745 1.355 1.005 ;
        RECT 1.130 0.730 1.300 0.745 ;
        POLYGON 1.130 0.730 1.230 0.730 1.230 0.630 ;
        RECT 1.230 0.000 1.300 0.730 ;
      LAYER via ;
        RECT 1.170 0.745 1.355 1.005 ;
      LAYER met2 ;
        RECT 0.000 1.005 1.300 1.030 ;
        RECT -0.055 0.745 1.355 1.005 ;
        RECT 0.000 0.580 1.300 0.745 ;
    END
  END VPWR
  OBS
      LAYER met2 ;
        RECT 0.000 1.600 1.300 2.055 ;
  END
END sky130_fd_bd_sram__sram_sp_colenda_cent
END LIBRARY

