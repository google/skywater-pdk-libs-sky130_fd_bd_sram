magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1271 1882 1587
<< psubdiffcont >>
rect 460 299 494 316
<< polycont >>
rect 567 262 601 292
<< locali >>
rect 594 174 611 175
rect 594 141 611 142
use sky130_fd_bd_sram__sram_dp_swldrv_mcon  sky130_fd_bd_sram__sram_dp_swldrv_mcon_0
timestamp 0
transform 1 0 216 0 1 14
box -9 -4 223 268
use sky130_fd_bd_sram__sram_dp_mcon_05  sky130_fd_bd_sram__sram_dp_mcon_05_0
timestamp 0
transform 0 1 0 -1 0 259
box -17 0 17 17
use sky130_fd_bd_sram__sram_dp_swldrv_strap2  sky130_fd_bd_sram__sram_dp_swldrv_strap2_0
timestamp 0
transform 1 0 0 0 1 0
box 0 0 74 316
use sky130_fd_bd_sram__sram_dp_swldrv_p1m_siz  sky130_fd_bd_sram__sram_dp_swldrv_p1m_siz_0
timestamp 0
transform 1 0 611 0 1 0
box -52 24 -33 293
use sky130_fd_bd_sram__sram_dp_swldrv_p1lic  sky130_fd_bd_sram__sram_dp_swldrv_p1lic_0
timestamp 0
transform 1 0 611 0 -1 316
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_p1m_ser  sky130_fd_bd_sram__sram_dp_swldrv_p1m_ser_0
timestamp 0
transform 1 0 611 0 1 -1
box -52 54 -34 293
use sky130_fd_bd_sram__sram_dp_swldrv_coreid  sky130_fd_bd_sram__sram_dp_swldrv_coreid_0
timestamp 0
transform 1 0 385 0 1 0
box 0 0 1 1
use sky130_fd_bd_sram__sram_dp_swldrv_met2_lwl  sky130_fd_bd_sram__sram_dp_swldrv_met2_lwl_0
timestamp 0
transform 1 0 611 0 -1 316
box -137 121 0 185
use sky130_fd_bd_sram__sram_dp_swldrv_base  sky130_fd_bd_sram__sram_dp_swldrv_base_0
timestamp 0
transform 1 0 611 0 1 0
box -611 0 0 316
use sky130_fd_bd_sram__sram_dp_swldrv_met23_2a  sky130_fd_bd_sram__sram_dp_swldrv_met23_2a_0
timestamp 0
transform 1 0 611 0 1 0
box -622 -11 11 327
use sky130_fd_bd_sram__sram_dp_swldrv_tap  sky130_fd_bd_sram__sram_dp_swldrv_tap_0
timestamp 0
transform 1 0 0 0 1 269
box 0 -62 519 47
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_swldrv_opt4a.gds
string GDS_END 10794
string GDS_START 10060
<< end >>
