magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1260 -1260 1884 1734
<< metal1 >>
rect 78 0 114 474
rect 150 0 186 474
rect 222 300 258 474
rect 214 256 266 300
rect 214 158 266 204
rect 222 0 258 158
rect 294 0 330 474
rect 366 0 402 474
<< via1 >>
rect 214 204 266 256
<< metal2 >>
rect 0 256 624 284
rect 0 204 214 256
rect 266 204 624 256
rect 0 174 624 204
<< labels >>
flabel metal1 s 78 196 114 244 0 FreeSans 2000 0 0 0 BL0
port 0 nsew
flabel metal1 s 294 196 330 244 0 FreeSans 2000 0 0 0 BL1
port 1 nsew
flabel metal1 s 150 196 186 244 0 FreeSans 2000 0 0 0 BR0
port 2 nsew
flabel metal1 s 366 196 402 244 0 FreeSans 2000 0 0 0 BR1
port 3 nsew
flabel metal2 s 311 214 342 248 0 FreeSans 2000 0 0 0 VDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 624 474
string GDS_FILE sky130_fd_bd_sram__openram_dp_cell_cap_col.gds
string GDS_END 1816
string GDS_START 174
<< end >>
