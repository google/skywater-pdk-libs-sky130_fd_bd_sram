magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1230 -1321 2792 1792
<< nwell >>
rect 622 -60 1532 532
<< pwell >>
rect 270 -17 352 19
<< nmos >>
rect 406 273 554 303
rect 406 201 554 231
rect 406 129 554 159
rect 406 57 554 87
<< pmos >>
rect 792 233 1016 263
rect 1166 233 1390 263
rect 792 145 1016 175
rect 1166 145 1390 175
<< ndiff >>
rect 406 351 554 359
rect 406 317 467 351
rect 501 317 554 351
rect 406 303 554 317
rect 406 231 554 273
rect 406 159 554 201
rect 406 87 554 129
rect 406 17 554 57
rect 406 -17 469 17
rect 503 -17 554 17
rect 406 -51 554 -17
<< pdiff >>
rect 792 315 1016 323
rect 792 281 887 315
rect 921 281 1016 315
rect 792 263 1016 281
rect 1166 315 1390 323
rect 1166 281 1261 315
rect 1295 281 1390 315
rect 1166 263 1390 281
rect 792 221 1016 233
rect 792 187 887 221
rect 921 187 1016 221
rect 792 175 1016 187
rect 1166 220 1390 233
rect 1166 186 1261 220
rect 1295 186 1390 220
rect 1166 175 1390 186
rect 792 129 1016 145
rect 792 95 887 129
rect 921 95 1016 129
rect 792 87 1016 95
rect 1166 133 1390 145
rect 1166 99 1261 133
rect 1295 99 1390 133
rect 1166 91 1390 99
<< ndiffc >>
rect 467 317 501 351
rect 469 -17 503 17
<< pdiffc >>
rect 887 281 921 315
rect 1261 281 1295 315
rect 887 187 921 221
rect 1261 186 1295 220
rect 887 95 921 129
rect 1261 99 1295 133
<< psubdiff >>
rect 270 17 352 19
rect 270 -17 294 17
rect 328 -17 352 17
rect 1238 17 1320 19
rect 1238 0 1262 17
rect 1296 0 1320 17
<< nsubdiff >>
rect 1238 -17 1262 0
rect 1296 -17 1320 0
rect 1238 -21 1320 -17
<< psubdiffcont >>
rect 294 -17 328 17
<< nsubdiffcont >>
rect 1262 -17 1296 17
<< poly >>
rect 324 323 378 339
rect 324 289 334 323
rect 368 303 378 323
rect 603 338 1121 368
rect 603 303 633 338
rect 368 289 406 303
rect 324 273 406 289
rect 554 273 633 303
rect 228 251 282 267
rect 228 217 238 251
rect 272 231 282 251
rect 1091 263 1121 338
rect 674 233 792 263
rect 1016 233 1042 263
rect 1091 234 1166 263
rect 1092 233 1166 234
rect 1390 233 1416 263
rect 674 231 704 233
rect 272 217 406 231
rect 228 201 406 217
rect 554 201 704 231
rect 132 179 186 195
rect 132 145 142 179
rect 176 159 186 179
rect 1090 175 1142 176
rect 738 159 792 175
rect 176 145 406 159
rect 132 129 406 145
rect 554 145 792 159
rect 1016 145 1042 175
rect 1090 145 1166 175
rect 1390 145 1416 175
rect 554 129 766 145
rect 36 107 90 123
rect 36 73 46 107
rect 80 87 90 107
rect 1090 144 1142 145
rect 80 73 406 87
rect 36 57 406 73
rect 554 71 676 87
rect 1090 72 1120 144
rect 1070 71 1122 72
rect 554 57 1122 71
rect 646 41 1122 57
rect 1070 40 1122 41
<< polycont >>
rect 334 289 368 323
rect 238 217 272 251
rect 142 145 176 179
rect 46 73 80 107
<< locali >>
rect 420 351 632 352
rect 318 289 334 323
rect 368 289 384 323
rect 420 317 467 351
rect 501 317 632 351
rect 592 315 632 317
rect 592 281 887 315
rect 921 281 1040 315
rect 1182 281 1261 315
rect 1295 281 1472 315
rect 222 217 238 251
rect 272 217 288 251
rect 719 192 753 281
rect 719 190 754 192
rect 126 145 142 179
rect 176 145 192 179
rect 715 128 754 190
rect 870 187 887 221
rect 921 187 937 221
rect 1244 220 1311 221
rect 1244 186 1261 220
rect 1295 186 1311 220
rect 1244 185 1311 186
rect 1244 132 1261 133
rect 870 128 887 129
rect 30 73 46 107
rect 80 73 96 107
rect 715 95 887 128
rect 921 95 938 129
rect 1182 99 1261 132
rect 1295 99 1312 133
rect 1182 98 1269 99
rect 715 94 895 95
rect 270 17 550 20
rect 270 -17 294 17
rect 328 -17 462 17
rect 503 -17 550 17
rect 270 -18 550 -17
rect 1260 17 1296 33
rect 1260 -17 1262 17
rect 1260 -33 1296 -17
<< viali >>
rect 887 187 921 221
rect 1261 186 1295 220
rect 462 -17 469 17
rect 469 -17 496 17
rect 1262 -17 1296 17
<< metal1 >>
rect 454 17 504 359
rect 454 -17 462 17
rect 496 -17 504 17
rect 454 -61 504 -17
rect 880 221 928 353
rect 880 187 887 221
rect 921 187 928 221
rect 880 -33 928 187
rect 1254 220 1302 363
rect 1254 186 1261 220
rect 1295 186 1302 220
rect 1254 17 1302 186
rect 1254 -17 1262 17
rect 1296 -17 1302 17
rect 1254 -33 1302 -17
<< labels >>
rlabel metal1 s 462 -51 498 -35 4 GND
port 4 nsew
rlabel metal1 s 902 -11 902 -11 4 VDD
port 5 nsew
rlabel metal1 s 1278 57 1278 57 4 VDD
port 5 nsew
rlabel locali s 350 305 350 305 4 A
port 0 nsew
rlabel locali s 254 233 254 233 4 B
port 1 nsew
rlabel locali s 158 161 158 161 4 C
port 2 nsew
rlabel locali s 64 89 64 89 4 D
port 3 nsew
rlabel locali s 1442 298 1442 298 4 Z
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 1522 395
string GDS_FILE sky130_fd_bd_sram__openram_dp_nand4_dec.gds
string GDS_END 6436
string GDS_START 170
<< end >>
