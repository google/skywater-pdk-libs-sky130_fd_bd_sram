magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1271 -1271 1500 1645
<< via1 >>
rect -11 -11 26 26
<< metal2 >>
rect 0 294 240 385
rect 0 26 240 217
rect 26 0 240 26
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_colend_half_met23_optb.gds
string GDS_END 386
string GDS_START 190
<< end >>
