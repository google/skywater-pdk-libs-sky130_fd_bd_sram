# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_colend_half_optb
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_colend_half_optb ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  1.310000 BY  1.925000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.585000 0.420000 1.925000 ;
      RECT 0.070000 0.000000 0.590000 0.095000 ;
      RECT 0.210000 0.345000 0.380000 0.515000 ;
      RECT 0.730000 0.000000 1.200000 0.095000 ;
      RECT 0.840000 0.585000 1.200000 1.925000 ;
      RECT 1.115000 0.515000 1.200000 0.585000 ;
    LAYER mcon ;
      RECT 0.000000 0.775000 0.085000 0.945000 ;
      RECT 0.395000 0.000000 0.565000 0.085000 ;
      RECT 0.755000 0.000000 0.925000 0.085000 ;
      RECT 1.115000 1.645000 1.200000 1.815000 ;
    LAYER met1 ;
      RECT -0.055000 0.730000 0.130000 0.990000 ;
      RECT  0.395000 0.000000 0.565000 0.085000 ;
      RECT  0.755000 0.000000 0.925000 0.085000 ;
      RECT  1.070000 1.565000 1.255000 1.825000 ;
    LAYER met2 ;
      RECT -0.055000 0.730000 0.130000 0.990000 ;
      RECT  1.070000 1.565000 1.255000 1.825000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 1.200000 0.205000 ;
    LAYER nwell ;
      RECT 0.720000 0.000000 1.200000 1.345000 ;
    LAYER pwell ;
      RECT 0.000000 0.715000 0.400000 1.505000 ;
      RECT 0.000000 1.505000 1.200000 1.795000 ;
      RECT 0.190000 0.585000 0.400000 0.715000 ;
  END
END sky130_fd_bd_sram__sram_dp_colend_half_optb
END LIBRARY
