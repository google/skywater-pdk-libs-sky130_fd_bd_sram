# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_rowend
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_rowend ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  1.355000 BY  1.580000 ;
  PIN vpwr
    ANTENNADIFFAREA  0.021600 ;
    PORT
      LAYER met2 ;
        RECT -0.055000 1.025000 1.300000 1.285000 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0.000000 0.705000 0.085000 0.875000 ;
      RECT 0.305000 0.605000 0.475000 0.775000 ;
      RECT 0.305000 0.965000 0.475000 1.135000 ;
      RECT 0.395000 0.200000 0.905000 0.370000 ;
      RECT 0.565000 0.620000 0.735000 0.790000 ;
      RECT 0.565000 0.960000 0.735000 1.130000 ;
    LAYER mcon ;
      RECT 0.565000 0.200000 0.735000 0.370000 ;
    LAYER met1 ;
      POLYGON  0.270000 0.600000 0.270000 0.540000 0.210000 0.540000 ;
      POLYGON  0.380000 0.600000 0.500000 0.600000 0.380000 0.480000 ;
      POLYGON  0.500000 0.610000 0.510000 0.610000 0.500000 0.600000 ;
      POLYGON  0.520000 0.100000 0.550000 0.100000 0.550000 0.070000 ;
      POLYGON  0.540000 0.440000 0.540000 0.420000 0.520000 0.420000 ;
      POLYGON  0.750000 0.100000 0.780000 0.100000 0.750000 0.070000 ;
      POLYGON  0.760000 0.440000 0.780000 0.420000 0.760000 0.420000 ;
      POLYGON  0.790000 0.610000 0.800000 0.610000 0.800000 0.600000 ;
      POLYGON  0.800000 0.600000 0.920000 0.600000 0.920000 0.480000 ;
      POLYGON  1.030000 0.600000 1.090000 0.540000 1.030000 0.540000 ;
      RECT -0.055000 1.025000 0.130000 1.285000 ;
      RECT  0.000000 0.000000 0.070000 0.635000 ;
      RECT  0.000000 0.635000 0.105000 0.990000 ;
      RECT  0.000000 0.990000 0.130000 1.025000 ;
      RECT  0.000000 1.285000 0.130000 1.315000 ;
      RECT  0.000000 1.315000 0.070000 1.580000 ;
      RECT  0.210000 0.000000 0.380000 0.540000 ;
      RECT  0.270000 0.540000 0.380000 0.600000 ;
      RECT  0.270000 0.600000 0.500000 0.610000 ;
      RECT  0.270000 0.610000 0.510000 1.580000 ;
      RECT  0.520000 0.100000 0.780000 0.420000 ;
      RECT  0.540000 0.420000 0.760000 0.440000 ;
      RECT  0.550000 0.070000 0.750000 0.100000 ;
      RECT  0.790000 0.610000 1.030000 1.580000 ;
      RECT  0.800000 0.600000 1.030000 0.610000 ;
      RECT  0.920000 0.000000 1.090000 0.540000 ;
      RECT  0.920000 0.540000 1.030000 0.600000 ;
    LAYER met2 ;
      RECT 0.000000 0.295000 1.300000 0.465000 ;
      RECT 0.000000 0.635000 1.300000 0.855000 ;
      RECT 0.520000 0.120000 0.780000 0.295000 ;
    LAYER nwell ;
      RECT 0.000000 0.000000 1.300000 1.580000 ;
    LAYER via ;
      RECT 0.520000 0.150000 0.780000 0.410000 ;
  END
END sky130_fd_bd_sram__sram_sp_rowend
END LIBRARY
