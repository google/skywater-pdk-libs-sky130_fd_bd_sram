* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_sram_dff CLK D Q Q_N
X0 a_547_102# a_28_102# gnd gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X1 a_239_76# CLK gnd gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X2 vdd a_47_611# a_28_102# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X3 gnd a_28_102# a_389_102# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X4 gnd Q a_739_102# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X5 Q Q_N gnd gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X6 a_389_712# a_239_76# a_47_611# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X7 a_47_611# a_239_76# a_197_102# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X8 Q_N CLK a_547_102# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X9 a_739_102# a_239_76# Q_N gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X10 a_547_712# a_28_102# vdd vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X11 a_239_76# CLK vdd vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X12 a_197_102# D gnd gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X13 vdd a_28_102# a_389_712# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X14 vdd Q a_739_712# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X15 gnd a_47_611# a_28_102# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X16 Q Q_N vdd vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X17 Q_N a_239_76# a_547_712# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X18 a_47_611# CLK a_197_712# vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X19 a_739_712# CLK Q_N vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X20 a_389_102# CLK a_47_611# gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X21 a_197_712# D vdd vdd sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
.ends
