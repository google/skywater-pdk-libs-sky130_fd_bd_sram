
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_sense_amp" ******************************

.SUBCKT sky130_fd_bd_sram__openram_sense_amp bl br dout en vdd gnd
X1000 gnd en a_56_432# gnd sky130_fd_pr__nfet_01v8 W=0.65u L=0.15u m=1
X1001 a_56_432# dint_bar dint gnd sky130_fd_pr__nfet_01v8 W=0.65u L=0.15u m=1
X1002 dint_bar dint a_56_432# gnd sky130_fd_pr__nfet_01v8 W=0.65u L=0.15u m=1

X1003 vdd dint_bar dint vdd sky130_fd_pr__pfet_01v8 W=1.26u L=0.15u m=1
X1004 dint_bar dint vdd vdd sky130_fd_pr__pfet_01v8 W=1.26u L=0.15u m=1

X1005 bl en dint vdd sky130_fd_pr__pfet_01v8 W=2u L=0.15u m=1
X1006 dint_bar en br vdd sky130_fd_pr__pfet_01v8 W=2u L=0.15u m=1

X1007 vdd dint_bar dout vdd sky130_fd_pr__pfet_01v8 W=1.26u L=0.15u m=1
X1008 dout dint_bar gnd gnd sky130_fd_pr__nfet_01v8 W=0.65u L=0.15u m=1

.ENDS sky130_fd_bd_sram__openram_sense_amp
