# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_nand3_dec
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_nand3_dec ;
  ORIGIN  0.360000 -0.175000 ;
  SIZE  6.965000 BY  1.580000 ;
  PIN GND
    ANTENNADIFFAREA  0.374750 ;
    PORT
      LAYER met1 ;
        RECT 0.890000 -0.220000 1.120000 1.840000 ;
      LAYER pwell ;
        RECT -0.320000 1.300000 -0.050000 1.715000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.844200 ;
    PORT
      LAYER met1 ;
        RECT 3.360000 0.070000 3.600000 1.840000 ;
        RECT 5.520000 0.070000 5.760000 1.840000 ;
      LAYER nwell ;
        RECT 2.070000 -0.300000 6.610000 2.370000 ;
    END
  END VDD
  OBS
    LAYER li1 ;
      RECT -0.350000 0.880000 -0.020000 1.050000 ;
      RECT -0.270000 1.300000 -0.100000 1.670000 ;
      RECT -0.270000 1.670000  0.900000 1.840000 ;
      RECT  0.200000 0.430000  0.530000 0.600000 ;
      RECT  0.200000 1.330000  0.530000 1.500000 ;
      RECT  0.700000 1.455000  1.360000 1.650000 ;
      RECT  0.700000 1.650000  0.900000 1.670000 ;
      RECT  0.710000 0.305000  6.610000 0.475000 ;
      RECT  1.630000 1.215000  1.970000 1.300000 ;
      RECT  1.630000 1.300000  2.055000 1.510000 ;
      RECT  2.555000 0.475000  2.725000 1.275000 ;
      RECT  2.555000 1.275000  3.650000 1.440000 ;
      RECT  2.555000 1.440000  3.435000 1.445000 ;
      RECT  3.310000 0.770000  5.805000 0.940000 ;
      RECT  3.310000 1.270000  3.650000 1.275000 ;
      RECT  4.610000 1.215000  4.950000 1.300000 ;
      RECT  4.610000 1.300000  5.035000 1.510000 ;
      RECT  5.550000 1.360000  5.740000 1.690000 ;
    LAYER mcon ;
      RECT 0.920000 1.465000 1.090000 1.635000 ;
      RECT 1.710000 1.275000 1.880000 1.445000 ;
      RECT 3.395000 0.770000 3.565000 0.940000 ;
      RECT 4.690000 1.275000 4.860000 1.445000 ;
      RECT 5.555000 0.770000 5.725000 0.940000 ;
      RECT 5.555000 1.440000 5.725000 1.610000 ;
    LAYER met1 ;
      RECT 1.630000 1.135000 1.975000 1.450000 ;
      RECT 1.630000 1.450000 1.970000 1.510000 ;
      RECT 4.610000 1.135000 4.955000 1.450000 ;
      RECT 4.610000 1.450000 4.950000 1.510000 ;
    LAYER met2 ;
      RECT 1.630000 1.135000 1.975000 1.300000 ;
      RECT 1.630000 1.300000 5.045000 1.440000 ;
      RECT 4.610000 1.135000 4.955000 1.300000 ;
    LAYER via ;
      RECT 1.670000 1.170000 1.930000 1.430000 ;
      RECT 4.650000 1.170000 4.910000 1.430000 ;
  END
END sky130_fd_bd_sram__openram_nand3_dec
END LIBRARY
