# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_corner_met2
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_corner_met2 ;
  ORIGIN  0.055000 -0.020000 ;
  SIZE  1.355000 BY  2.035000 ;
  OBS
    LAYER met1 ;
      RECT -0.055000 0.745000 0.130000 1.005000 ;
      RECT  0.270000 1.200000 0.530000 1.460000 ;
      RECT  0.800000 0.120000 1.060000 0.380000 ;
    LAYER met2 ;
      RECT -0.055000 0.745000 1.300000 1.005000 ;
      RECT  0.000000 0.020000 1.300000 0.405000 ;
      RECT  0.000000 0.580000 1.300000 0.745000 ;
      RECT  0.000000 1.005000 1.300000 1.030000 ;
      RECT  0.000000 1.180000 1.300000 1.460000 ;
      RECT  0.000000 1.600000 1.300000 2.055000 ;
  END
END sky130_fd_bd_sram__sram_sp_corner_met2
END LIBRARY
