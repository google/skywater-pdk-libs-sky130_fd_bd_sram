* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__sram_dp_blkinv_base m1_0_0# a_48_42# a_100_0# SUBS m1_298_0#
+ a_100_72# a_100_158# a_559_24#
X0 a_419_146# a_48_42# a_100_72# SUBS sky130_fd_pr__nfet_01v8 w=310000u l=150000u
X1 a_100_72# a_48_42# a_419_0# SUBS sky130_fd_pr__nfet_01v8 w=310000u l=150000u
X2 a_100_158# a_48_42# a_100_72# w_0_0# sky130_fd_pr__pfet_01v8 w=930000u l=150000u
X3 a_100_72# a_48_42# a_100_0# w_0_0# sky130_fd_pr__pfet_01v8 w=930000u l=150000u
.ends
* Top level circuit sky130_fd_bd_sram__sram_dp_blkinv_opt2a
Xsky130_fd_bd_sram__sram_dp_blkinv_base_0 sky130_fd_bd_sram__sram_dp_blkinv_base_0/m1_0_0#
+ sky130_fd_bd_sram__sram_dp_blkinv_base_0/a_48_42# li_210_n3# SUBS sky130_fd_bd_sram__sram_dp_blkinv_base_0/m1_298_0#
+ sky130_fd_bd_sram__sram_dp_blkinv_base_0/m1_298_0# a_100_158# sky130_fd_bd_sram__sram_dp_blkinv_base_0/a_559_24#
+ sky130_fd_bd_sram__sram_dp_blkinv_base
.end
