* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_bd_sram__openram_sense_amp BL BR DOUT EN GND VDD
X0 GND a_154_1298# DOUT GND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_154_1298# a_96_1689# VDD VDD sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X2 BL EN a_96_1689# VDD sky130_fd_pr__pfet_01v8 w=2e+06u l=150000u
X3 GND EN a_184_1689# GND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_184_1689# a_154_1298# a_96_1689# GND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_154_1298# EN BR VDD sky130_fd_pr__pfet_01v8 w=2e+06u l=150000u
X6 a_154_1298# a_96_1689# a_184_1689# GND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VDD a_154_1298# a_96_1689# VDD sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X8 VDD a_154_1298# DOUT VDD sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
.ends
