
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_sense_amp" ******************************

.SUBCKT sky130_fd_bd_sram__openram_sense_amp bl br dout en vdd gnd
M1000 gnd en a_56_432# gnd nshort W=0.65 L=0.15 m=1 mult=1
M1001 a_56_432# dint_bar dint gnd nshort W=0.65 L=0.15 m=1 mult=1
M1002 dint_bar dint a_56_432# gnd nshort W=0.65 L=0.15 m=1 mult=1

M1003 vdd dint_bar dint vdd pshort W=1.26 L=0.15 m=1 mult=1
M1004 dint_bar dint vdd vdd pshort W=1.26 L=0.15 m=1 mult=1

M1005 bl en dint vdd pshort W=2 L=0.15 m=1 mult=1
M1006 dint_bar en br vdd pshort W=2 L=0.15 m=1 mult=1

M1007 vdd dint_bar dout vdd pshort W=1.26 L=0.15 m=1 mult=1
M1008 dout dint_bar gnd gnd nshort W=0.65 L=0.15 m=1 mult=1

.ENDS sky130_fd_bd_sram__openram_sense_amp
