# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cell_opt1
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cell_opt1 ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  1.310000 BY  1.580000 ;
  PIN bl
    ANTENNADIFFAREA  0.016800 ;
    PORT
      LAYER met1 ;
        RECT 0.300000 1.435000 0.540000 1.580000 ;
        RECT 0.350000 0.000000 0.490000 1.435000 ;
    END
  END bl
  PIN br
    ANTENNADIFFAREA  0.016800 ;
    PORT
      LAYER met1 ;
        RECT 0.660000 0.000000 0.900000 0.145000 ;
        RECT 0.710000 0.145000 0.850000 1.580000 ;
    END
  END br
  PIN vgnd
    ANTENNADIFFAREA  0.080800 ;
    PORT
      LAYER met2 ;
        RECT -0.055000 0.635000 1.200000 0.855000 ;
        RECT -0.055000 0.855000 0.290000 0.895000 ;
    END
  END vgnd
  PIN vnb
    PORT
      LAYER pwell ;
        RECT 0.010000 0.170000 0.060000 0.230000 ;
    END
  END vnb
  PIN vpb
    PORT
      LAYER nwell ;
        RECT 0.690000 0.065000 1.200000 1.515000 ;
        RECT 0.720000 0.000000 1.200000 0.065000 ;
        RECT 0.720000 1.515000 1.200000 1.580000 ;
    END
  END vpb
  PIN vpwr
    ANTENNADIFFAREA  0.064000 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1.065000 1.255000 1.285000 ;
        RECT 0.955000 1.025000 1.255000 1.065000 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0.000000 0.705000 0.085000 0.875000 ;
      RECT 0.190000 0.000000 0.330000 0.085000 ;
      RECT 0.190000 0.310000 0.330000 0.395000 ;
      RECT 0.190000 0.395000 0.355000 0.480000 ;
      RECT 0.190000 1.100000 0.355000 1.185000 ;
      RECT 0.190000 1.185000 0.330000 1.270000 ;
      RECT 0.190000 1.495000 0.330000 1.580000 ;
      RECT 0.335000 1.495000 0.505000 1.580000 ;
      RECT 0.535000 0.520000 0.705000 0.670000 ;
      RECT 0.535000 0.910000 0.705000 1.060000 ;
      RECT 0.695000 0.000000 0.865000 0.085000 ;
      RECT 0.870000 0.305000 1.010000 0.475000 ;
      RECT 0.870000 1.105000 1.010000 1.275000 ;
      RECT 1.115000 0.705000 1.200000 0.875000 ;
    LAYER met1 ;
      POLYGON  1.085000 0.645000 1.095000 0.645000 1.095000 0.635000 ;
      RECT -0.055000 0.635000 0.130000 0.895000 ;
      RECT  0.000000 0.000000 0.070000 0.605000 ;
      RECT  0.000000 0.605000 0.130000 0.635000 ;
      RECT  0.000000 0.895000 0.130000 0.925000 ;
      RECT  0.000000 0.925000 0.070000 1.580000 ;
      RECT  1.070000 0.990000 1.200000 1.025000 ;
      RECT  1.070000 1.025000 1.255000 1.285000 ;
      RECT  1.070000 1.285000 1.200000 1.315000 ;
      RECT  1.085000 0.645000 1.200000 0.990000 ;
      RECT  1.095000 0.635000 1.200000 0.645000 ;
      RECT  1.130000 0.000000 1.200000 0.635000 ;
      RECT  1.130000 1.315000 1.200000 1.580000 ;
    LAYER met2 ;
      RECT 0.000000 0.295000 1.200000 0.465000 ;
  END
END sky130_fd_bd_sram__sram_sp_cell_opt1
END LIBRARY
