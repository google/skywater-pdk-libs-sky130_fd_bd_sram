# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_cell_1rw_1r
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_cell_1rw_1r ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.120000 BY  1.975000 ;
  OBS
    LAYER li1 ;
      RECT -0.085000 -0.085000 0.085000 0.085000 ;
      RECT -0.085000  1.100000 0.085000 1.270000 ;
      RECT  0.210000 -0.085000 0.380000 0.085000 ;
      RECT  0.210000  0.320000 0.380000 0.470000 ;
      RECT  0.210000  0.705000 0.380000 0.875000 ;
      RECT  0.210000  1.495000 0.380000 1.665000 ;
      RECT  0.210000  1.890000 0.380000 1.975000 ;
      RECT  0.395000  1.890000 0.565000 2.060000 ;
      RECT  0.535000  1.035000 0.695000 1.065000 ;
      RECT  0.545000  1.065000 0.695000 1.205000 ;
      RECT  0.755000  1.890000 0.925000 2.060000 ;
      RECT  0.980000  0.695000 1.120000 0.865000 ;
      RECT  0.980000  1.100000 1.285000 1.270000 ;
      RECT  0.980000  1.505000 1.120000 1.675000 ;
      RECT  1.390000  1.120000 1.525000 1.290000 ;
      RECT  1.475000  0.310000 1.645000 0.480000 ;
      RECT  1.705000  1.165000 1.855000 1.305000 ;
      RECT  1.705000  1.305000 1.865000 1.335000 ;
      RECT  1.835000  0.310000 2.005000 0.480000 ;
      RECT  2.020000 -0.085000 2.190000 0.085000 ;
      RECT  2.020000  0.310000 2.190000 0.480000 ;
      RECT  2.020000  0.705000 2.190000 0.875000 ;
      RECT  2.020000  1.495000 2.190000 1.665000 ;
      RECT  2.020000  1.900000 2.190000 1.975000 ;
      RECT  2.315000 -0.085000 2.485000 0.085000 ;
      RECT  2.330000  1.105000 2.485000 1.265000 ;
      RECT  2.470000  0.590000 2.740000 0.715000 ;
      RECT  2.470000  0.715000 2.640000 0.760000 ;
      RECT  2.470000  1.610000 2.640000 1.655000 ;
      RECT  2.470000  1.655000 2.740000 1.780000 ;
      RECT  2.570000 -0.085000 2.740000 0.085000 ;
      RECT  2.570000  0.545000 2.740000 0.590000 ;
      RECT  2.570000  1.780000 2.740000 1.825000 ;
      RECT  2.825000 -0.085000 2.995000 0.085000 ;
      RECT  2.825000  1.105000 3.015000 1.265000 ;
      RECT  2.845000  1.100000 3.015000 1.105000 ;
      RECT  2.845000  1.265000 3.015000 1.270000 ;
    LAYER mcon ;
      RECT 1.115000 1.100000 1.285000 1.270000 ;
      RECT 2.470000 0.590000 2.640000 0.760000 ;
    LAYER met1 ;
      POLYGON  2.575000  0.895000 2.655000  0.815000 2.575000 0.815000 ;
      POLYGON  2.575000  1.555000 2.655000  1.555000 2.575000 1.475000 ;
      RECT -0.210000 -0.520000 0.210000  2.100000 ;
      RECT  0.390000 -0.520000 0.570000  2.100000 ;
      RECT  0.750000 -0.520000 0.930000  2.100000 ;
      RECT  1.110000 -0.520000 1.290000  2.100000 ;
      RECT  1.470000 -0.520000 1.650000  2.100000 ;
      RECT  1.830000 -0.520000 2.010000  2.100000 ;
      RECT  2.190000 -0.190000 3.120000  0.190000 ;
      RECT  2.190000  0.485000 2.655000  0.815000 ;
      RECT  2.190000  0.815000 2.575000  0.895000 ;
      RECT  2.190000  1.475000 2.575000  1.555000 ;
      RECT  2.190000  1.555000 2.655000  1.885000 ;
      RECT  2.750000  0.980000 3.120000  1.390000 ;
      RECT  2.835000 -0.520000 3.120000 -0.190000 ;
      RECT  2.835000  0.190000 3.120000  0.980000 ;
      RECT  2.835000  1.390000 3.120000  2.100000 ;
    LAYER met2 ;
      RECT -0.210000 -0.275000 3.120000 0.275000 ;
      RECT -0.210000  0.515000 3.120000 0.755000 ;
      RECT -0.210000  0.995000 2.020000 1.065000 ;
      RECT -0.210000  1.065000 3.120000 1.305000 ;
      RECT -0.210000  1.305000 2.020000 1.375000 ;
      RECT -0.210000  1.615000 3.120000 1.855000 ;
      RECT  2.190000  0.755000 2.600000 0.825000 ;
      RECT  2.190000  1.545000 2.600000 1.615000 ;
      RECT  2.770000  0.995000 3.120000 1.065000 ;
      RECT  2.770000  1.305000 3.120000 1.375000 ;
    LAYER nwell ;
      RECT 0.720000 -0.395000 1.680000 1.975000 ;
    LAYER pwell ;
      RECT 0.190000 -0.195000 0.400000 0.195000 ;
    LAYER pwell ;
      RECT 2.000000 -0.195000 2.210000 0.195000 ;
    LAYER via ;
      RECT -0.130000 -0.130000 0.130000 0.130000 ;
      RECT -0.130000  1.055000 0.130000 1.315000 ;
      RECT  2.265000  0.540000 2.525000 0.800000 ;
      RECT  2.265000  1.570000 2.525000 1.830000 ;
      RECT  2.270000 -0.130000 2.530000 0.130000 ;
      RECT  2.780000 -0.130000 3.040000 0.130000 ;
      RECT  2.805000  1.055000 3.065000 1.315000 ;
  END
END sky130_fd_bd_sram__openram_cell_1rw_1r
END LIBRARY
