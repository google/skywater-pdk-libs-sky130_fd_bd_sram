
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_nand3_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_nand3_dec
.subckt sky130_fd_bd_sram__openram_nand3_dec A B C Z vdd gnd

X1001 Z A a_n346_328# gnd sky130_fd_pr__nfet_01v8 W=0.74u L=0.15u m=1
X1002 a_n346_256# C gnd gnd sky130_fd_pr__nfet_01v8 W=0.74u L=0.15u m=1
X1003 a_n346_328# B a_n346_256# gnd sky130_fd_pr__nfet_01v8 W=0.74u L=0.15u m=1
X1000 Z B vdd vdd sky130_fd_pr__pfet_01v8 W=1.12u L=0.15u m=1
X1004 Z A vdd vdd sky130_fd_pr__pfet_01v8 W=1.12u L=0.15u m=1
X1005 Z C vdd vdd sky130_fd_pr__pfet_01v8 W=1.12u L=0.15u m=1
.ends

