# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_cornera
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_cornera ;
  ORIGIN  0.055000  0.000000 ;
  SIZE  1.355000 BY  2.055000 ;
  PIN vnb
    PORT
      LAYER met2 ;
        RECT 0.000000 0.020000 1.300000 0.405000 ;
    END
  END vnb
  PIN vpb
    ANTENNADIFFAREA  0.414475 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1.180000 1.300000 1.460000 ;
      LAYER nwell ;
        RECT 0.000000 0.000000 0.445000 2.055000 ;
    END
  END vpb
  PIN vpwr
    PORT
      LAYER met2 ;
        RECT -0.055000 0.745000 1.300000 1.005000 ;
        RECT  0.000000 0.580000 1.300000 0.745000 ;
        RECT  0.000000 1.005000 1.300000 1.030000 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0.000000 0.275000 1.130000 0.810000 ;
      RECT 0.000000 0.990000 0.340000 1.160000 ;
      RECT 0.000000 1.160000 1.300000 1.875000 ;
      RECT 0.160000 0.000000 1.130000 0.275000 ;
      RECT 0.520000 0.810000 1.130000 0.990000 ;
    LAYER mcon ;
      RECT 0.285000 1.250000 0.455000 1.420000 ;
      RECT 0.285000 1.610000 0.455000 1.780000 ;
      RECT 0.790000 0.755000 0.960000 0.925000 ;
      RECT 0.900000 0.055000 1.070000 0.225000 ;
    LAYER met1 ;
      POLYGON  0.070000 0.730000 0.170000 0.730000 0.070000 0.630000 ;
      POLYGON  0.090000 1.105000 0.170000 1.025000 0.090000 1.025000 ;
      POLYGON  0.250000 1.205000 0.255000 1.205000 0.255000 1.200000 ;
      POLYGON  0.255000 1.200000 0.310000 1.200000 0.310000 1.145000 ;
      POLYGON  0.310000 0.495000 0.310000 0.395000 0.210000 0.395000 ;
      POLYGON  0.380000 0.170000 0.550000 0.170000 0.380000 0.000000 ;
      POLYGON  0.760000 0.160000 0.800000 0.160000 0.800000 0.120000 ;
      POLYGON  0.800000 0.120000 0.865000 0.120000 0.865000 0.055000 ;
      POLYGON  0.865000 0.055000 0.920000 0.055000 0.920000 0.000000 ;
      POLYGON  0.990000 0.465000 1.075000 0.380000 0.990000 0.380000 ;
      POLYGON  0.990000 1.215000 1.060000 1.215000 0.990000 1.145000 ;
      POLYGON  1.075000 0.380000 1.090000 0.365000 1.075000 0.365000 ;
      RECT -0.055000 0.745000 0.170000 1.005000 ;
      RECT  0.000000 0.000000 0.070000 0.730000 ;
      RECT  0.000000 0.730000 0.170000 0.745000 ;
      RECT  0.000000 1.005000 0.170000 1.025000 ;
      RECT  0.000000 1.025000 0.090000 2.055000 ;
      RECT  0.210000 0.000000 0.380000 0.170000 ;
      RECT  0.210000 0.170000 0.550000 0.395000 ;
      RECT  0.250000 1.205000 0.550000 2.055000 ;
      RECT  0.255000 1.200000 0.550000 1.205000 ;
      RECT  0.310000 0.395000 0.550000 1.200000 ;
      RECT  0.760000 0.160000 1.090000 0.365000 ;
      RECT  0.760000 0.365000 1.075000 0.380000 ;
      RECT  0.760000 0.380000 0.990000 1.215000 ;
      RECT  0.760000 1.215000 1.060000 2.055000 ;
      RECT  0.800000 0.120000 1.090000 0.160000 ;
      RECT  0.865000 0.055000 1.090000 0.120000 ;
      RECT  0.920000 0.000000 1.090000 0.055000 ;
    LAYER met2 ;
      RECT 0.000000 1.600000 1.300000 2.055000 ;
    LAYER via ;
      RECT 0.270000 1.200000 0.530000 1.460000 ;
      RECT 0.800000 0.120000 1.060000 0.380000 ;
  END
END sky130_fd_bd_sram__sram_sp_cornera
END LIBRARY
