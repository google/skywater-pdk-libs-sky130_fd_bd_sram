* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_cent_m2.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_cent_m2
.ends
