# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_dp_nand2_dec
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_dp_nand2_dec ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.380000 BY  1.975000 ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.350000 1.410000 0.680000 1.580000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.350000 0.870000 0.680000 1.040000 ;
    END
  END B
  PIN GND
    ANTENNADIFFAREA  0.393800 ;
    PORT
      LAYER met1 ;
        RECT 1.230000 -0.150000 1.470000 2.010000 ;
      LAYER pwell ;
        RECT 1.140000 -0.090000 1.560000 0.090000 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA  0.415800 ;
    PORT
      LAYER met1 ;
        RECT 3.350000 -0.160000 3.600000 2.010000 ;
      LAYER nwell ;
        RECT 2.060000 -0.280000 4.440000 2.380000 ;
    END
  END VDD
  PIN Z
    ANTENNADIFFAREA  0.826800 ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.570000 4.440000 1.740000 ;
        RECT 2.545000 0.670000 2.860000 0.675000 ;
        RECT 2.545000 0.675000 3.425000 0.680000 ;
        RECT 2.545000 0.680000 3.640000 0.845000 ;
        RECT 2.545000 0.845000 2.990000 0.850000 ;
        RECT 2.545000 0.850000 2.715000 1.570000 ;
        RECT 3.300000 0.845000 3.640000 0.850000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT 1.040000  0.710000 1.700000 0.880000 ;
      RECT 1.180000 -0.090000 1.560000 0.090000 ;
      RECT 3.300000 -0.095000 3.650000 0.095000 ;
      RECT 3.300000  1.130000 3.635000 1.300000 ;
    LAYER mcon ;
      RECT 1.265000 -0.085000 1.435000 0.085000 ;
      RECT 1.270000  0.710000 1.440000 0.880000 ;
      RECT 3.385000  1.130000 3.555000 1.300000 ;
      RECT 3.395000 -0.085000 3.565000 0.085000 ;
  END
END sky130_fd_bd_sram__openram_dp_nand2_dec
END LIBRARY
