VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__openram_sp_cell_p1_serifs
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__openram_sp_cell_p1_serifs ;
  ORIGIN -0.010 -0.125 ;
  SIZE 0.965 BY 0.395 ;
END sky130_fd_bd_sram__openram_sp_cell_p1_serifs
END LIBRARY

