magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -1735 -1320 2725 1735
<< nwell >>
rect 1086 474 1465 475
rect 414 -60 1465 474
<< pwell >>
rect -59 260 -5 343
<< nmos >>
rect 128 250 276 280
rect -384 158 -232 188
rect 128 178 276 208
rect 128 106 276 136
<< pmos >>
rect 584 206 808 236
rect 1050 205 1275 238
rect 584 106 808 136
rect 1050 106 1275 136
<< ndiff >>
rect 128 327 276 351
rect -384 237 -232 261
rect 128 293 191 327
rect 225 293 276 327
rect 128 280 276 293
rect -384 203 -323 237
rect -289 203 -232 237
rect -384 188 -232 203
rect 128 208 276 250
rect -384 142 -232 158
rect -384 108 -326 142
rect -292 108 -232 142
rect 128 136 276 178
rect -384 98 -232 108
rect 128 95 276 106
rect 128 61 189 95
rect 223 61 276 95
rect 128 53 276 61
<< pdiff >>
rect 584 288 808 296
rect 584 254 679 288
rect 713 254 808 288
rect 584 236 808 254
rect 1050 285 1275 296
rect 1050 251 1145 285
rect 1179 251 1275 285
rect 1050 238 1275 251
rect 584 188 808 206
rect 584 154 679 188
rect 713 154 808 188
rect 584 136 808 154
rect 1050 188 1275 205
rect 1050 154 1145 188
rect 1179 154 1275 188
rect 1050 136 1275 154
rect 584 95 808 106
rect 584 61 679 95
rect 713 61 808 95
rect 584 46 808 61
rect 1050 95 1275 106
rect 1050 61 1145 95
rect 1179 61 1275 95
rect 1050 46 1275 61
<< ndiffc >>
rect 191 293 225 327
rect -323 203 -289 237
rect -326 108 -292 142
rect 189 61 223 95
<< pdiffc >>
rect 679 254 713 288
rect 1145 251 1179 285
rect 679 154 713 188
rect 1145 154 1179 188
rect 679 61 713 95
rect 1145 61 1179 95
<< psubdiff >>
rect -59 318 -5 343
rect -59 284 -49 318
rect -15 284 -5 318
rect -59 260 -5 284
<< nsubdiff >>
rect 1380 318 1414 351
rect 1380 258 1414 284
<< psubdiffcont >>
rect -49 284 -15 318
<< nsubdiffcont >>
rect 1380 284 1414 318
<< poly >>
rect 46 300 100 316
rect 46 266 56 300
rect 90 280 100 300
rect 331 300 386 316
rect 331 280 342 300
rect 90 266 128 280
rect 46 250 128 266
rect 276 266 342 280
rect 376 266 386 300
rect 928 300 982 316
rect 276 250 386 266
rect -469 190 -415 206
rect -469 156 -459 190
rect -425 188 -415 190
rect -194 230 -139 246
rect -194 196 -183 230
rect -149 197 -139 230
rect -64 210 -10 226
rect -149 196 -138 197
rect -194 188 -138 196
rect -425 158 -384 188
rect -232 158 -138 188
rect -64 176 -54 210
rect -20 208 -10 210
rect 928 266 938 300
rect 972 266 982 300
rect 470 208 584 236
rect -20 178 128 208
rect 276 206 584 208
rect 808 206 834 236
rect 928 234 982 266
rect 276 178 500 206
rect -20 176 -10 178
rect -64 160 -10 176
rect -425 156 -415 158
rect -469 140 -415 156
rect 940 136 970 234
rect 1024 205 1050 238
rect 1275 205 1395 238
rect 1341 200 1395 205
rect 1341 166 1351 200
rect 1385 166 1395 200
rect 1341 150 1395 166
rect 46 120 128 136
rect 46 86 56 120
rect 90 106 128 120
rect 276 106 584 136
rect 808 106 834 136
rect 940 106 1050 136
rect 1275 106 1301 136
rect 90 86 100 106
rect 46 70 100 86
<< polycont >>
rect 56 266 90 300
rect 342 266 376 300
rect -459 156 -425 190
rect -183 196 -149 230
rect -54 176 -20 210
rect 938 266 972 300
rect 1351 166 1385 200
rect 56 86 90 120
<< locali >>
rect -337 318 1 351
rect -337 316 -49 318
rect -337 240 -290 316
rect -59 284 -49 316
rect -15 284 1 318
rect 140 327 272 330
rect -59 268 1 284
rect 40 266 56 300
rect 90 266 106 300
rect 140 293 191 327
rect 225 293 272 327
rect 140 291 272 293
rect 326 300 411 302
rect 326 255 342 300
rect 376 260 411 300
rect 922 300 1007 302
rect 511 288 687 289
rect 376 255 394 260
rect 326 243 394 255
rect 511 255 679 288
rect -374 237 -242 240
rect -374 203 -330 237
rect -289 203 -242 237
rect -374 201 -242 203
rect -199 230 -114 232
rect -475 156 -459 190
rect -425 156 -409 190
rect -199 185 -183 230
rect -149 190 -114 230
rect -149 185 -131 190
rect -199 173 -131 185
rect -70 176 -54 210
rect -20 176 -4 210
rect -373 142 -243 145
rect -373 108 -330 142
rect -292 108 -243 142
rect -373 106 -243 108
rect 40 86 56 120
rect 90 86 106 120
rect 511 95 545 255
rect 662 254 679 255
rect 713 254 730 288
rect 922 255 938 300
rect 972 260 1007 300
rect 972 255 990 260
rect 922 243 990 255
rect 1129 251 1145 285
rect 1179 251 1263 285
rect 1364 283 1380 318
rect 1414 283 1430 318
rect 1364 280 1430 283
rect 662 154 679 188
rect 713 154 1145 188
rect 1179 154 1195 188
rect 1229 95 1263 251
rect 1335 200 1403 202
rect 1335 155 1351 200
rect 1385 155 1403 200
rect 1335 143 1403 155
rect 142 61 189 95
rect 223 61 679 95
rect 713 61 1145 95
rect 1179 61 1356 95
<< viali >>
rect 191 293 225 327
rect 342 266 376 289
rect 342 255 376 266
rect -330 203 -323 237
rect -323 203 -296 237
rect -183 196 -149 219
rect -183 185 -149 196
rect -330 108 -326 142
rect -326 108 -296 142
rect 938 266 972 289
rect 938 255 972 266
rect 1380 284 1414 317
rect 1380 283 1414 284
rect 679 154 713 188
rect 1145 154 1179 188
rect 1351 166 1385 189
rect 1351 155 1385 166
<< metal1 >>
rect 179 327 237 340
rect 179 293 191 327
rect 225 293 237 327
rect -337 237 -290 293
rect -337 203 -330 237
rect -296 203 -290 237
rect -337 185 -290 203
rect -199 220 -131 232
rect -199 219 -130 220
rect -199 216 -183 219
rect -149 216 -130 219
rect -199 164 -191 216
rect -139 164 -130 216
rect -199 157 -130 164
rect -343 142 -250 151
rect -343 108 -330 142
rect -296 128 -250 142
rect 179 128 237 293
rect 326 290 394 302
rect 326 289 395 290
rect 326 286 342 289
rect 376 286 395 289
rect 326 234 334 286
rect 386 234 395 286
rect 326 227 395 234
rect 672 188 720 368
rect 1138 324 1186 349
rect 1138 317 1460 324
rect 922 290 990 302
rect 922 289 991 290
rect 922 286 938 289
rect 972 286 991 289
rect 922 234 930 286
rect 982 234 991 286
rect 922 227 991 234
rect 1138 283 1380 317
rect 1414 283 1460 317
rect 1138 276 1460 283
rect 672 154 679 188
rect 713 154 720 188
rect -296 108 277 128
rect -343 100 277 108
rect 672 14 720 154
rect 1138 188 1186 276
rect 1138 154 1145 188
rect 1179 154 1186 188
rect 1138 14 1186 154
rect 1335 189 1403 202
rect 1335 186 1351 189
rect 1385 186 1403 189
rect 1335 134 1343 186
rect 1395 134 1403 186
rect 1335 127 1403 134
<< via1 >>
rect -191 185 -183 216
rect -183 185 -149 216
rect -149 185 -139 216
rect -191 164 -139 185
rect 334 255 342 286
rect 342 255 376 286
rect 376 255 386 286
rect 334 234 386 255
rect 930 255 938 286
rect 938 255 972 286
rect 972 255 982 286
rect 930 234 982 255
rect 1343 155 1351 186
rect 1351 155 1385 186
rect 1385 155 1395 186
rect 1343 134 1395 155
<< metal2 >>
rect 326 286 1009 288
rect 326 234 334 286
rect 386 260 930 286
rect 386 234 395 260
rect 326 227 395 234
rect 922 234 930 260
rect 982 260 1009 286
rect 982 234 991 260
rect 922 227 991 234
rect -199 216 -130 218
rect -199 164 -191 216
rect -139 199 -130 216
rect -139 186 1403 199
rect -139 171 1343 186
rect -139 164 -130 171
rect -199 157 -130 164
rect 1335 134 1343 171
rect 1395 134 1403 186
rect 1335 127 1403 134
<< labels >>
rlabel corelocali s -445 176 -445 176 4 D
rlabel corelocali s 70 284 70 284 4 C
rlabel corelocali s -40 196 -40 196 4 B
rlabel corelocali s 70 106 70 106 4 A
rlabel corelocali s 1328 78 1328 78 4 Z
rlabel metal1 s 677 338 715 356 4 VDD
port 1 nsew
rlabel metal1 s 1430 281 1448 319 4 VDD
port 1 nsew
rlabel metal1 s -333 266 -295 284 4 GND
port 0 nsew
<< properties >>
string FIXED_BBOX -475 35 1460 351
string GDS_FILE sky130_fd_bd_sram__openram_nand4_dec.gds
string GDS_END 8988
string GDS_START 162
<< end >>
