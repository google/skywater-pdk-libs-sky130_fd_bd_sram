# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_wls_half
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_wls_half ;
  ORIGIN  0.035000  0.000000 ;
  SIZE  0.645000 BY  0.500000 ;
  OBS
    LAYER li1 ;
      RECT 0.170000 0.090000 0.540000 0.405000 ;
    LAYER mcon ;
      RECT 0.170000 0.195000 0.340000 0.365000 ;
    LAYER met1 ;
      POLYGON  0.275000 0.500000 0.355000 0.420000 0.275000 0.420000 ;
      RECT -0.035000 0.145000 0.355000 0.405000 ;
      RECT  0.100000 0.090000 0.355000 0.145000 ;
      RECT  0.100000 0.405000 0.355000 0.420000 ;
      RECT  0.100000 0.420000 0.275000 0.500000 ;
    LAYER met2 ;
      RECT -0.035000 0.145000 0.610000 0.360000 ;
      RECT -0.035000 0.360000 0.300000 0.405000 ;
      RECT  0.100000 0.120000 0.610000 0.145000 ;
      RECT  0.100000 0.405000 0.300000 0.430000 ;
    LAYER met3 ;
      RECT 0.100000 0.000000 0.610000 0.205000 ;
  END
END sky130_fd_bd_sram__sram_dp_wls_half
END LIBRARY
