* NGSPICE file created from sky130_fd_bd_sram__sram_sp_corner_ce.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_corner_ce
.ends
