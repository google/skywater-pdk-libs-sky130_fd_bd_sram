# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_sp_colend_cent_ce
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_sp_colend_cent_ce ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.300000 BY  2.055000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.275000 1.300000 0.810000 ;
      RECT 0.000000 0.990000 1.300000 1.875000 ;
      RECT 0.135000 0.015000 1.200000 0.275000 ;
    LAYER mcon ;
      RECT 0.295000 1.345000 0.465000 1.515000 ;
      RECT 0.295000 1.705000 0.465000 1.875000 ;
      RECT 0.790000 0.280000 0.960000 0.450000 ;
      RECT 0.790000 0.640000 0.960000 0.810000 ;
    LAYER met1 ;
      POLYGON 0.070000 0.730000 0.170000 0.730000 0.070000 0.630000 ;
      POLYGON 0.090000 1.100000 0.170000 1.020000 0.090000 1.020000 ;
      POLYGON 0.250000 1.155000 0.305000 1.155000 0.305000 1.100000 ;
      POLYGON 0.305000 1.100000 0.310000 1.100000 0.310000 1.095000 ;
      POLYGON 0.310000 0.480000 0.310000 0.380000 0.210000 0.380000 ;
      POLYGON 0.380000 0.170000 0.550000 0.170000 0.380000 0.000000 ;
      POLYGON 0.750000 0.170000 0.920000 0.170000 0.920000 0.000000 ;
      POLYGON 0.990000 0.480000 1.090000 0.380000 0.990000 0.380000 ;
      POLYGON 0.990000 1.155000 1.050000 1.155000 0.990000 1.095000 ;
      POLYGON 1.130000 0.730000 1.230000 0.730000 1.230000 0.630000 ;
      POLYGON 1.200000 1.095000 1.200000 1.025000 1.130000 1.025000 ;
      POLYGON 1.210000 1.105000 1.210000 1.095000 1.200000 1.095000 ;
      RECT 0.000000 0.000000 0.070000 0.730000 ;
      RECT 0.000000 0.730000 0.170000 1.020000 ;
      RECT 0.000000 1.020000 0.090000 2.055000 ;
      RECT 0.210000 0.000000 0.380000 0.170000 ;
      RECT 0.210000 0.170000 0.550000 0.380000 ;
      RECT 0.250000 1.155000 0.550000 2.055000 ;
      RECT 0.305000 1.100000 0.550000 1.155000 ;
      RECT 0.310000 0.380000 0.550000 1.100000 ;
      RECT 0.750000 0.170000 1.090000 0.380000 ;
      RECT 0.750000 0.380000 0.990000 1.155000 ;
      RECT 0.750000 1.155000 1.050000 2.055000 ;
      RECT 0.920000 0.000000 1.090000 0.170000 ;
      RECT 1.130000 0.730000 1.300000 1.025000 ;
      RECT 1.200000 1.025000 1.300000 1.095000 ;
      RECT 1.210000 1.095000 1.300000 2.055000 ;
      RECT 1.230000 0.000000 1.300000 0.730000 ;
    LAYER nwell ;
      RECT 0.000000 0.000000 1.300000 2.055000 ;
  END
END sky130_fd_bd_sram__sram_sp_colend_cent_ce
END LIBRARY
