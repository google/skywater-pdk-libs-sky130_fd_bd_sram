
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_nand2_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_nand2_dec
.subckt sky130_fd_bd_sram__openram_nand2_dec A B Z vdd gnd

M1001 Z B vdd vdd pshort W=1.12 L=0.15 m=1 mult=1
M1002 vdd A Z vdd pshort W=1.12 L=0.15 m=1 mult=1
M1000 Z A a_n722_276# gnd nshort W=0.74 L=0.15 m=1 mult=1
M1003 a_n722_276# B gnd gnd nshort W=0.74 L=0.15 m=1 mult=1
.ends

