# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_cell_opt5
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_cell_opt5 ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  2.510000 BY  1.690000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.625000 0.070000 0.705000 ;
      RECT 0.000000 0.705000 0.085000 0.875000 ;
      RECT 0.000000 0.875000 0.070000 0.955000 ;
      RECT 0.070000 0.000000 0.590000 0.125000 ;
      RECT 0.070000 0.295000 1.865000 0.470000 ;
      RECT 0.070000 1.505000 1.670000 1.580000 ;
      RECT 0.210000 0.470000 1.865000 0.475000 ;
      RECT 0.210000 0.475000 0.380000 1.365000 ;
      RECT 0.210000 1.495000 0.380000 1.505000 ;
      RECT 0.490000 1.455000 1.670000 1.505000 ;
      RECT 0.535000 0.670000 0.705000 1.105000 ;
      RECT 0.535000 1.105000 2.190000 1.110000 ;
      RECT 0.535000 1.110000 2.330000 1.285000 ;
      RECT 0.730000 0.000000 2.330000 0.075000 ;
      RECT 0.730000 0.075000 1.910000 0.125000 ;
      RECT 0.860000 0.655000 1.540000 0.925000 ;
      RECT 1.695000 0.475000 1.865000 0.910000 ;
      RECT 1.810000 1.455000 2.330000 1.580000 ;
      RECT 2.020000 0.075000 2.190000 0.085000 ;
      RECT 2.020000 0.215000 2.190000 1.105000 ;
      RECT 2.315000 0.705000 2.400000 0.875000 ;
      RECT 2.330000 0.215000 2.400000 0.705000 ;
      RECT 2.330000 0.875000 2.400000 0.970000 ;
    LAYER mcon ;
      RECT 0.395000 0.000000 0.565000 0.085000 ;
      RECT 0.755000 0.000000 0.925000 0.085000 ;
      RECT 1.115000 0.705000 1.285000 0.875000 ;
      RECT 1.475000 1.495000 1.645000 1.580000 ;
      RECT 1.835000 1.495000 2.005000 1.580000 ;
    LAYER met1 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.210000 0.130000 ;
      RECT -0.055000  1.450000 0.210000 1.580000 ;
      RECT -0.055000  1.580000 0.130000 1.635000 ;
      RECT  0.000000  0.130000 0.210000 1.450000 ;
      RECT  0.390000  0.000000 0.570000 1.580000 ;
      RECT  0.750000  0.000000 0.930000 1.580000 ;
      RECT  1.110000  0.000000 1.290000 1.580000 ;
      RECT  1.470000  0.000000 1.650000 1.580000 ;
      RECT  1.830000  0.000000 2.010000 1.580000 ;
      RECT  2.190000  0.000000 2.400000 0.660000 ;
      RECT  2.190000  0.660000 2.455000 0.920000 ;
      RECT  2.190000  0.920000 2.400000 1.580000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.205000 0.130000 ;
      RECT -0.055000  1.450000 1.860000 1.580000 ;
      RECT -0.055000  1.580000 0.130000 1.635000 ;
      RECT  0.000000  0.130000 0.205000 0.185000 ;
      RECT  0.000000  0.605000 0.780000 0.845000 ;
      RECT  0.000000  1.395000 1.860000 1.450000 ;
      RECT  0.540000  0.120000 2.400000 0.360000 ;
      RECT  0.540000  0.360000 0.780000 0.605000 ;
      RECT  1.620000  0.740000 2.455000 0.920000 ;
      RECT  1.620000  0.920000 2.400000 0.980000 ;
      RECT  1.620000  0.980000 1.860000 1.395000 ;
      RECT  2.195000  0.600000 2.400000 0.660000 ;
      RECT  2.195000  0.660000 2.455000 0.740000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 2.400000 0.205000 ;
      RECT 0.000000 0.505000 2.400000 1.075000 ;
      RECT 0.000000 1.375000 2.400000 1.580000 ;
    LAYER nwell ;
      RECT 0.720000 0.000000 1.680000 1.580000 ;
    LAYER via ;
      RECT 2.270000 0.660000 2.455000 0.920000 ;
  END
END sky130_fd_bd_sram__sram_dp_cell_opt5
END LIBRARY
