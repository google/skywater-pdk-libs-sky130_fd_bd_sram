magic
tech sky130A
magscale 1 2
timestamp 1621288236
<< dnwell >>
rect 0 0 260 411
<< nwell >>
rect 0 0 89 411
<< nsubdiff >>
rect 0 368 59 375
rect 0 334 17 368
rect 51 334 59 368
rect 0 300 59 334
rect 0 266 17 300
rect 51 266 59 300
rect 0 232 59 266
rect 0 198 17 232
rect 51 198 59 232
rect 0 94 59 198
<< nsubdiffcont >>
rect 17 334 51 368
rect 17 266 51 300
rect 17 198 51 232
<< poly >>
rect 16 68 150 84
rect 16 54 32 68
rect 0 34 32 54
rect 66 34 100 68
rect 134 34 150 68
rect 0 24 150 34
rect 16 18 150 24
<< polycont >>
rect 32 34 66 68
rect 100 34 134 68
<< locali >>
rect 0 368 260 375
rect 0 334 17 368
rect 51 356 260 368
rect 51 334 57 356
rect 0 322 57 334
rect 91 322 260 356
rect 0 300 260 322
rect 0 266 17 300
rect 51 284 260 300
rect 51 266 57 284
rect 0 250 57 266
rect 91 250 260 284
rect 0 232 260 250
rect 0 198 17 232
rect 51 198 68 232
rect 104 185 226 198
rect 104 162 158 185
rect 0 151 158 162
rect 192 151 226 185
rect 0 68 226 151
rect 0 55 32 68
rect 66 34 100 68
rect 134 45 226 68
rect 134 34 180 45
rect 32 11 180 34
rect 214 11 226 45
rect 32 0 226 11
<< viali >>
rect 57 322 91 356
rect 57 250 91 284
rect 158 151 192 185
rect 180 11 214 45
<< metal1 >>
rect 0 205 18 411
rect 50 356 110 411
rect 50 322 57 356
rect 91 322 110 356
rect 50 291 110 322
rect 50 241 55 291
rect 105 241 110 291
tri 50 229 62 241 ne
tri 18 205 34 221 sw
rect 0 200 34 205
rect 25 150 34 200
rect 0 146 34 150
rect 0 0 14 146
tri 14 126 34 146 nw
tri 42 79 62 99 se
rect 62 79 110 241
rect 42 34 110 79
rect 42 0 76 34
tri 76 0 110 34 nw
rect 152 243 212 411
rect 152 185 198 243
tri 198 229 212 243 nw
rect 152 151 158 185
rect 192 151 198 185
rect 152 75 198 151
tri 198 75 216 93 sw
rect 152 32 161 75
rect 211 73 216 75
tri 216 73 218 75 sw
rect 211 45 218 73
tri 152 25 159 32 ne
rect 159 25 161 32
tri 159 11 173 25 ne
rect 173 11 180 25
rect 214 11 218 45
tri 173 0 184 11 ne
rect 184 0 218 11
<< via1 >>
rect 55 284 105 291
rect 55 250 57 284
rect 57 250 91 284
rect 91 250 105 284
rect 55 241 105 250
rect -10 150 25 200
rect 161 45 211 75
rect 161 25 180 45
rect 180 25 211 45
<< metal2 >>
rect 0 320 260 411
rect 0 291 260 292
rect 0 241 55 291
rect 105 241 260 291
rect 0 236 260 241
rect 0 200 260 206
rect 25 150 260 200
rect 0 116 260 150
rect 0 75 260 81
rect 0 25 161 75
rect 211 25 260 75
rect 0 4 260 25
<< labels >>
rlabel metal1 s 0 0 14 19 4 VPWR
rlabel metal1 s 50 375 110 411 4 VPB
rlabel metal1 s 152 375 212 411 4 VNB
<< end >>
