# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_bd_sram__sram_dp_colend_opt6
  CLASS BLOCK ;
  FOREIGN sky130_fd_bd_sram__sram_dp_colend_opt6 ;
  ORIGIN  0.055000  0.055000 ;
  SIZE  2.510000 BY  1.980000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.585000 0.420000 1.925000 ;
      RECT 0.070000 0.000000 1.670000 0.095000 ;
      RECT 0.210000 0.345000 0.380000 0.515000 ;
      RECT 0.840000 0.585000 1.560000 1.925000 ;
      RECT 1.115000 0.515000 1.285000 0.585000 ;
      RECT 1.810000 0.000000 2.330000 0.095000 ;
      RECT 1.980000 0.585000 2.400000 1.925000 ;
      RECT 2.020000 0.345000 2.190000 0.515000 ;
    LAYER mcon ;
      RECT 0.000000 0.775000 0.085000 0.945000 ;
      RECT 1.115000 1.645000 1.285000 1.815000 ;
      RECT 1.475000 0.000000 1.645000 0.085000 ;
      RECT 1.835000 0.000000 2.005000 0.085000 ;
      RECT 2.315000 0.775000 2.400000 0.945000 ;
    LAYER met1 ;
      POLYGON  0.090000  1.150000 0.210000 1.030000 0.090000 1.030000 ;
      POLYGON  0.270000  1.225000 0.345000 1.225000 0.345000 1.150000 ;
      POLYGON  0.345000  1.150000 0.390000 1.150000 0.390000 1.105000 ;
      POLYGON  0.450000  1.300000 0.570000 1.180000 0.450000 1.180000 ;
      POLYGON  0.630000  1.375000 0.705000 1.375000 0.705000 1.300000 ;
      POLYGON  0.705000  1.300000 0.750000 1.300000 0.750000 1.255000 ;
      POLYGON  0.810000  1.450000 0.930000 1.330000 0.810000 1.330000 ;
      POLYGON  0.990000  1.525000 1.065000 1.525000 1.065000 1.450000 ;
      POLYGON  1.065000  1.450000 1.110000 1.450000 1.110000 1.405000 ;
      POLYGON  1.290000  1.525000 1.410000 1.525000 1.290000 1.405000 ;
      POLYGON  1.545000  1.405000 1.545000 1.330000 1.470000 1.330000 ;
      POLYGON  1.590000  1.450000 1.590000 1.405000 1.545000 1.405000 ;
      POLYGON  1.650000  1.375000 1.770000 1.375000 1.650000 1.255000 ;
      POLYGON  1.905000  1.255000 1.905000 1.180000 1.830000 1.180000 ;
      POLYGON  1.950000  1.300000 1.950000 1.255000 1.905000 1.255000 ;
      POLYGON  2.010000  1.225000 2.130000 1.225000 2.010000 1.105000 ;
      POLYGON  2.265000  1.105000 2.265000 1.030000 2.190000 1.030000 ;
      POLYGON  2.310000  1.150000 2.310000 1.105000 2.265000 1.105000 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.210000 0.130000 ;
      RECT -0.055000  0.730000 0.210000 0.990000 ;
      RECT  0.000000  0.130000 0.210000 0.730000 ;
      RECT  0.000000  0.990000 0.210000 1.030000 ;
      RECT  0.000000  1.030000 0.090000 1.925000 ;
      RECT  0.270000  1.225000 0.450000 1.925000 ;
      RECT  0.345000  1.150000 0.570000 1.180000 ;
      RECT  0.345000  1.180000 0.450000 1.225000 ;
      RECT  0.390000  0.000000 0.570000 1.150000 ;
      RECT  0.630000  1.375000 0.810000 1.925000 ;
      RECT  0.705000  1.300000 0.930000 1.330000 ;
      RECT  0.705000  1.330000 0.810000 1.375000 ;
      RECT  0.750000  0.000000 0.930000 1.300000 ;
      RECT  0.990000  1.525000 1.410000 1.925000 ;
      RECT  1.065000  1.450000 1.290000 1.525000 ;
      RECT  1.110000  0.000000 1.290000 1.450000 ;
      RECT  1.470000  0.000000 1.650000 1.330000 ;
      RECT  1.545000  1.330000 1.650000 1.375000 ;
      RECT  1.545000  1.375000 1.770000 1.405000 ;
      RECT  1.590000  1.405000 1.770000 1.925000 ;
      RECT  1.830000  0.000000 2.010000 1.180000 ;
      RECT  1.905000  1.180000 2.010000 1.225000 ;
      RECT  1.905000  1.225000 2.130000 1.255000 ;
      RECT  1.950000  1.255000 2.130000 1.925000 ;
      RECT  2.190000  0.000000 2.400000 0.730000 ;
      RECT  2.190000  0.730000 2.455000 0.990000 ;
      RECT  2.190000  0.990000 2.400000 1.030000 ;
      RECT  2.265000  1.030000 2.400000 1.105000 ;
      RECT  2.310000  1.105000 2.400000 1.925000 ;
    LAYER met2 ;
      RECT -0.055000 -0.055000 0.130000 0.000000 ;
      RECT -0.055000  0.000000 0.205000 0.120000 ;
      RECT -0.055000  0.120000 2.400000 0.130000 ;
      RECT -0.055000  0.730000 2.455000 0.990000 ;
      RECT  0.000000  0.130000 2.400000 0.730000 ;
      RECT  0.000000  0.990000 2.400000 1.085000 ;
      RECT  0.000000  1.470000 2.400000 1.925000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 2.400000 0.205000 ;
    LAYER nwell ;
      RECT 0.720000 0.000000 1.680000 1.345000 ;
    LAYER pwell ;
      RECT 0.000000 0.715000 0.400000 1.505000 ;
      RECT 0.000000 1.505000 2.400000 1.795000 ;
      RECT 0.190000 0.585000 0.400000 0.715000 ;
    LAYER pwell ;
      RECT 2.000000 0.585000 2.210000 0.715000 ;
      RECT 2.000000 0.715000 2.400000 1.505000 ;
    LAYER via ;
      RECT 1.070000 1.565000 1.330000 1.825000 ;
      RECT 2.270000 0.730000 2.455000 0.990000 ;
  END
END sky130_fd_bd_sram__sram_dp_colend_opt6
END LIBRARY
