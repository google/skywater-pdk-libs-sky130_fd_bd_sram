magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -965 -1260 1661 1277
<< viali >>
rect 295 0 329 17
rect 367 0 401 17
<< properties >>
string GDS_FILE sky130_fd_bd_sram__sram_dp_horstrap_mcon.gds
string GDS_END 302
string GDS_START 170
<< end >>
